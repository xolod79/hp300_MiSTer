library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity videorom is
	generic(
		addr_width : integer := 8192;
		addr_bits  : integer := 13;
		data_width : integer := 8
        );
port(
    clk_i  : in std_logic;
    addr_i : in std_logic_vector(addr_bits-1 downto 0);
    data_o : out std_logic_vector(data_width-1 downto 0)
);
end videorom;

architecture rtl of videorom is

type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);
signal rom_i : rom_type := (
		x"39", -- 0
		x"00", -- 1
		x"04", -- 2
		x"00", -- 3
		x"04", -- 4
		x"00", -- 5
		x"04", -- 6
		x"00", -- 7
		x"03", -- 8
		x"00", -- 9
		x"02", -- a
		x"00", -- b
		x"01", -- c
		x"01", -- d
		x"01", -- e
		x"40", -- f
		x"00", -- 10
		x"01", -- 11
		x"01", -- 12
		x"00", -- 13
		x"00", -- 14
		x"00", -- 15
		x"00", -- 16
		x"00", -- 17
		x"00", -- 18
		x"00", -- 19
		x"00", -- 1a
		x"40", -- 1b
		x"00", -- 1c
		x"02", -- 1d
		x"01", -- 1e
		x"00", -- 1f
		x"00", -- 20
		x"00", -- 21
		x"00", -- 22
		x"00", -- 23
		x"00", -- 24
		x"00", -- 25
		x"00", -- 26
		x"00", -- 27
		x"00", -- 28
		x"00", -- 29
		x"00", -- 2a
		x"00", -- 2b
		x"00", -- 2c
		x"00", -- 2d
		x"00", -- 2e
		x"ff", -- 2f
		x"00", -- 30
		x"00", -- 31
		x"00", -- 32
		x"00", -- 33
		x"00", -- 34
		x"00", -- 35
		x"00", -- 36
		x"00", -- 37
		x"00", -- 38
		x"00", -- 39
		x"00", -- 3a
		x"00", -- 3b
		x"00", -- 3c
		x"00", -- 3d
		x"00", -- 3e
		x"00", -- 3f
		x"01", -- 40
		x"00", -- 41
		x"00", -- 42
		x"00", -- 43
		x"00", -- 44
		x"00", -- 45
		x"00", -- 46
		x"00", -- 47
		x"00", -- 48
		x"00", -- 49
		x"00", -- 4a
		x"00", -- 4b
		x"00", -- 4c
		x"00", -- 4d
		x"00", -- 4e
		x"00", -- 4f
		x"00", -- 50
		x"00", -- 51
		x"00", -- 52
		x"00", -- 53
		x"00", -- 54
		x"00", -- 55
		x"00", -- 56
		x"00", -- 57
		x"00", -- 58
		x"00", -- 59
		x"00", -- 5a
		x"00", -- 5b
		x"00", -- 5c
		x"00", -- 5d
		x"00", -- 5e
		x"00", -- 5f
		x"00", -- 60
		x"00", -- 61
		x"00", -- 62
		x"00", -- 63
		x"00", -- 64
		x"00", -- 65
		x"00", -- 66
		x"00", -- 67
		x"00", -- 68
		x"00", -- 69
		x"00", -- 6a
		x"00", -- 6b
		x"00", -- 6c
		x"00", -- 6d
		x"00", -- 6e
		x"00", -- 6f
		x"00", -- 70
		x"00", -- 71
		x"00", -- 72
		x"00", -- 73
		x"00", -- 74
		x"00", -- 75
		x"00", -- 76
		x"00", -- 77
		x"00", -- 78
		x"00", -- 79
		x"00", -- 7a
		x"00", -- 7b
		x"00", -- 7c
		x"00", -- 7d
		x"00", -- 7e
		x"20", -- 7f
		x"00", -- 80
		x"00", -- 81
		x"40", -- 82
		x"88", -- 83
		x"ff", -- 84
		x"00", -- 85
		x"00", -- 86
		x"00", -- 87
		x"40", -- 88
		x"8c", -- 89
		x"01", -- 8a
		x"00", -- 8b
		x"00", -- 8c
		x"00", -- 8d
		x"40", -- 8e
		x"90", -- 8f
		x"ff", -- 90
		x"00", -- 91
		x"00", -- 92
		x"00", -- 93
		x"40", -- 94
		x"ea", -- 95
		x"03", -- 96
		x"00", -- 97
		x"00", -- 98
		x"00", -- 99
		x"41", -- 9a
		x"42", -- 9b
		x"c0", -- 9c
		x"40", -- 9d
		x"00", -- 9e
		x"00", -- 9f
		x"41", -- a0
		x"46", -- a1
		x"90", -- a2
		x"05", -- a3
		x"00", -- a4
		x"00", -- a5
		x"41", -- a6
		x"4a", -- a7
		x"20", -- a8
		x"08", -- a9
		x"00", -- aa
		x"00", -- ab
		x"41", -- ac
		x"4e", -- ad
		x"70", -- ae
		x"07", -- af
		x"00", -- b0
		x"00", -- b1
		x"41", -- b2
		x"52", -- b3
		x"c3", -- b4
		x"00", -- b5
		x"00", -- b6
		x"00", -- b7
		x"41", -- b8
		x"56", -- b9
		x"90", -- ba
		x"03", -- bb
		x"00", -- bc
		x"00", -- bd
		x"41", -- be
		x"5a", -- bf
		x"20", -- c0
		x"04", -- c1
		x"00", -- c2
		x"00", -- c3
		x"41", -- c4
		x"5e", -- c5
		x"70", -- c6
		x"14", -- c7
		x"00", -- c8
		x"00", -- c9
		x"40", -- ca
		x"ac", -- cb
		x"00", -- cc
		x"00", -- cd
		x"00", -- ce
		x"00", -- cf
		x"40", -- d0
		x"84", -- d1
		x"01", -- d2
		x"00", -- d3
		x"80", -- d4
		x"00", -- d5
		x"40", -- d6
		x"80", -- d7
		x"ff", -- d8
		x"00", -- d9
		x"00", -- da
		x"00", -- db
		x"00", -- dc
		x"00", -- dd
		x"00", -- de
		x"00", -- df
		x"00", -- e0
		x"00", -- e1
		x"00", -- e2
		x"00", -- e3
		x"00", -- e4
		x"00", -- e5
		x"00", -- e6
		x"00", -- e7
		x"00", -- e8
		x"00", -- e9
		x"00", -- ea
		x"00", -- eb
		x"00", -- ec
		x"00", -- ed
		x"00", -- ee
		x"00", -- ef
		x"00", -- f0
		x"00", -- f1
		x"00", -- f2
		x"00", -- f3
		x"00", -- f4
		x"00", -- f5
		x"00", -- f6
		x"00", -- f7
		x"00", -- f8
		x"00", -- f9
		x"00", -- fa
		x"00", -- fb
		x"00", -- fc
		x"00", -- fd
		x"00", -- fe
		x"00", -- ff
		x"02", -- 100
		x"01", -- 101
		x"02", -- 102
		x"0f", -- 103
		x"02", -- 104
		x"22", -- 105
		x"19", -- 106
		x"10", -- 107
		x"08", -- 108
		x"01", -- 109
		x"00", -- 10a
		x"ff", -- 10b
		x"00", -- 10c
		x"48", -- 10d
		x"68", -- 10e
		x"58", -- 10f
		x"48", -- 110
		x"48", -- 111
		x"00", -- 112
		x"12", -- 113
		x"12", -- 114
		x"12", -- 115
		x"12", -- 116
		x"0c", -- 117
		x"00", -- 118
		x"00", -- 119
		x"00", -- 11a
		x"00", -- 11b
		x"00", -- 11c
		x"38", -- 11d
		x"40", -- 11e
		x"30", -- 11f
		x"08", -- 120
		x"70", -- 121
		x"00", -- 122
		x"12", -- 123
		x"12", -- 124
		x"1e", -- 125
		x"12", -- 126
		x"12", -- 127
		x"00", -- 128
		x"00", -- 129
		x"00", -- 12a
		x"00", -- 12b
		x"00", -- 12c
		x"38", -- 12d
		x"40", -- 12e
		x"30", -- 12f
		x"08", -- 130
		x"70", -- 131
		x"00", -- 132
		x"22", -- 133
		x"14", -- 134
		x"08", -- 135
		x"14", -- 136
		x"22", -- 137
		x"00", -- 138
		x"00", -- 139
		x"00", -- 13a
		x"00", -- 13b
		x"00", -- 13c
		x"78", -- 13d
		x"40", -- 13e
		x"70", -- 13f
		x"40", -- 140
		x"78", -- 141
		x"00", -- 142
		x"22", -- 143
		x"14", -- 144
		x"08", -- 145
		x"14", -- 146
		x"22", -- 147
		x"00", -- 148
		x"00", -- 149
		x"00", -- 14a
		x"00", -- 14b
		x"00", -- 14c
		x"78", -- 14d
		x"40", -- 14e
		x"70", -- 14f
		x"40", -- 150
		x"78", -- 151
		x"00", -- 152
		x"3e", -- 153
		x"08", -- 154
		x"08", -- 155
		x"08", -- 156
		x"08", -- 157
		x"00", -- 158
		x"00", -- 159
		x"00", -- 15a
		x"00", -- 15b
		x"00", -- 15c
		x"78", -- 15d
		x"40", -- 15e
		x"70", -- 15f
		x"40", -- 160
		x"78", -- 161
		x"00", -- 162
		x"1c", -- 163
		x"22", -- 164
		x"22", -- 165
		x"2a", -- 166
		x"1c", -- 167
		x"04", -- 168
		x"00", -- 169
		x"00", -- 16a
		x"00", -- 16b
		x"00", -- 16c
		x"30", -- 16d
		x"48", -- 16e
		x"78", -- 16f
		x"48", -- 170
		x"48", -- 171
		x"00", -- 172
		x"12", -- 173
		x"14", -- 174
		x"18", -- 175
		x"14", -- 176
		x"12", -- 177
		x"00", -- 178
		x"00", -- 179
		x"00", -- 17a
		x"00", -- 17b
		x"00", -- 17c
		x"00", -- 17d
		x"38", -- 17e
		x"44", -- 17f
		x"44", -- 180
		x"44", -- 181
		x"44", -- 182
		x"44", -- 183
		x"44", -- 184
		x"fe", -- 185
		x"10", -- 186
		x"00", -- 187
		x"00", -- 188
		x"00", -- 189
		x"00", -- 18a
		x"00", -- 18b
		x"00", -- 18c
		x"70", -- 18d
		x"48", -- 18e
		x"70", -- 18f
		x"48", -- 190
		x"70", -- 191
		x"00", -- 192
		x"0e", -- 193
		x"10", -- 194
		x"0c", -- 195
		x"02", -- 196
		x"1c", -- 197
		x"00", -- 198
		x"00", -- 199
		x"00", -- 19a
		x"00", -- 19b
		x"00", -- 19c
		x"48", -- 19d
		x"48", -- 19e
		x"78", -- 19f
		x"48", -- 1a0
		x"48", -- 1a1
		x"00", -- 1a2
		x"3e", -- 1a3
		x"08", -- 1a4
		x"08", -- 1a5
		x"08", -- 1a6
		x"08", -- 1a7
		x"00", -- 1a8
		x"00", -- 1a9
		x"00", -- 1aa
		x"00", -- 1ab
		x"00", -- 1ac
		x"40", -- 1ad
		x"40", -- 1ae
		x"40", -- 1af
		x"40", -- 1b0
		x"78", -- 1b1
		x"00", -- 1b2
		x"1e", -- 1b3
		x"10", -- 1b4
		x"1c", -- 1b5
		x"10", -- 1b6
		x"10", -- 1b7
		x"00", -- 1b8
		x"00", -- 1b9
		x"00", -- 1ba
		x"00", -- 1bb
		x"00", -- 1bc
		x"44", -- 1bd
		x"44", -- 1be
		x"28", -- 1bf
		x"28", -- 1c0
		x"10", -- 1c1
		x"00", -- 1c2
		x"3e", -- 1c3
		x"08", -- 1c4
		x"08", -- 1c5
		x"08", -- 1c6
		x"08", -- 1c7
		x"00", -- 1c8
		x"00", -- 1c9
		x"00", -- 1ca
		x"00", -- 1cb
		x"00", -- 1cc
		x"78", -- 1cd
		x"40", -- 1ce
		x"70", -- 1cf
		x"40", -- 1d0
		x"40", -- 1d1
		x"00", -- 1d2
		x"1e", -- 1d3
		x"10", -- 1d4
		x"1c", -- 1d5
		x"10", -- 1d6
		x"10", -- 1d7
		x"00", -- 1d8
		x"00", -- 1d9
		x"00", -- 1da
		x"00", -- 1db
		x"00", -- 1dc
		x"38", -- 1dd
		x"40", -- 1de
		x"40", -- 1df
		x"40", -- 1e0
		x"38", -- 1e1
		x"00", -- 1e2
		x"1c", -- 1e3
		x"12", -- 1e4
		x"1c", -- 1e5
		x"14", -- 1e6
		x"12", -- 1e7
		x"00", -- 1e8
		x"00", -- 1e9
		x"00", -- 1ea
		x"00", -- 1eb
		x"00", -- 1ec
		x"38", -- 1ed
		x"40", -- 1ee
		x"30", -- 1ef
		x"08", -- 1f0
		x"70", -- 1f1
		x"00", -- 1f2
		x"0c", -- 1f3
		x"12", -- 1f4
		x"12", -- 1f5
		x"12", -- 1f6
		x"0c", -- 1f7
		x"00", -- 1f8
		x"00", -- 1f9
		x"00", -- 1fa
		x"00", -- 1fb
		x"00", -- 1fc
		x"38", -- 1fd
		x"40", -- 1fe
		x"30", -- 1ff
		x"08", -- 200
		x"70", -- 201
		x"00", -- 202
		x"0e", -- 203
		x"04", -- 204
		x"04", -- 205
		x"04", -- 206
		x"0e", -- 207
		x"00", -- 208
		x"00", -- 209
		x"00", -- 20a
		x"00", -- 20b
		x"00", -- 20c
		x"70", -- 20d
		x"48", -- 20e
		x"48", -- 20f
		x"48", -- 210
		x"70", -- 211
		x"00", -- 212
		x"10", -- 213
		x"10", -- 214
		x"10", -- 215
		x"10", -- 216
		x"1e", -- 217
		x"00", -- 218
		x"00", -- 219
		x"00", -- 21a
		x"00", -- 21b
		x"00", -- 21c
		x"70", -- 21d
		x"48", -- 21e
		x"48", -- 21f
		x"48", -- 220
		x"70", -- 221
		x"00", -- 222
		x"04", -- 223
		x"0c", -- 224
		x"04", -- 225
		x"04", -- 226
		x"0e", -- 227
		x"00", -- 228
		x"00", -- 229
		x"00", -- 22a
		x"00", -- 22b
		x"00", -- 22c
		x"70", -- 22d
		x"48", -- 22e
		x"48", -- 22f
		x"48", -- 230
		x"70", -- 231
		x"0c", -- 232
		x"12", -- 233
		x"02", -- 234
		x"0c", -- 235
		x"10", -- 236
		x"1e", -- 237
		x"00", -- 238
		x"00", -- 239
		x"00", -- 23a
		x"00", -- 23b
		x"00", -- 23c
		x"70", -- 23d
		x"48", -- 23e
		x"48", -- 23f
		x"48", -- 240
		x"70", -- 241
		x"00", -- 242
		x"1c", -- 243
		x"02", -- 244
		x"0c", -- 245
		x"02", -- 246
		x"1c", -- 247
		x"00", -- 248
		x"00", -- 249
		x"00", -- 24a
		x"00", -- 24b
		x"00", -- 24c
		x"70", -- 24d
		x"48", -- 24e
		x"48", -- 24f
		x"48", -- 250
		x"70", -- 251
		x"00", -- 252
		x"14", -- 253
		x"14", -- 254
		x"1e", -- 255
		x"04", -- 256
		x"04", -- 257
		x"00", -- 258
		x"00", -- 259
		x"00", -- 25a
		x"00", -- 25b
		x"00", -- 25c
		x"48", -- 25d
		x"68", -- 25e
		x"58", -- 25f
		x"48", -- 260
		x"48", -- 261
		x"00", -- 262
		x"12", -- 263
		x"14", -- 264
		x"18", -- 265
		x"14", -- 266
		x"12", -- 267
		x"00", -- 268
		x"00", -- 269
		x"00", -- 26a
		x"00", -- 26b
		x"00", -- 26c
		x"38", -- 26d
		x"40", -- 26e
		x"30", -- 26f
		x"08", -- 270
		x"70", -- 271
		x"00", -- 272
		x"22", -- 273
		x"14", -- 274
		x"08", -- 275
		x"08", -- 276
		x"08", -- 277
		x"00", -- 278
		x"00", -- 279
		x"00", -- 27a
		x"00", -- 27b
		x"00", -- 27c
		x"78", -- 27d
		x"40", -- 27e
		x"70", -- 27f
		x"40", -- 280
		x"78", -- 281
		x"00", -- 282
		x"1c", -- 283
		x"12", -- 284
		x"1c", -- 285
		x"12", -- 286
		x"1c", -- 287
		x"00", -- 288
		x"00", -- 289
		x"00", -- 28a
		x"00", -- 28b
		x"00", -- 28c
		x"38", -- 28d
		x"40", -- 28e
		x"40", -- 28f
		x"40", -- 290
		x"38", -- 291
		x"00", -- 292
		x"12", -- 293
		x"1a", -- 294
		x"16", -- 295
		x"12", -- 296
		x"12", -- 297
		x"00", -- 298
		x"00", -- 299
		x"00", -- 29a
		x"00", -- 29b
		x"00", -- 29c
		x"78", -- 29d
		x"40", -- 29e
		x"70", -- 29f
		x"40", -- 2a0
		x"78", -- 2a1
		x"00", -- 2a2
		x"22", -- 2a3
		x"36", -- 2a4
		x"2a", -- 2a5
		x"22", -- 2a6
		x"22", -- 2a7
		x"00", -- 2a8
		x"00", -- 2a9
		x"00", -- 2aa
		x"00", -- 2ab
		x"00", -- 2ac
		x"38", -- 2ad
		x"40", -- 2ae
		x"30", -- 2af
		x"08", -- 2b0
		x"70", -- 2b1
		x"00", -- 2b2
		x"1c", -- 2b3
		x"12", -- 2b4
		x"1c", -- 2b5
		x"12", -- 2b6
		x"1c", -- 2b7
		x"00", -- 2b8
		x"00", -- 2b9
		x"00", -- 2ba
		x"00", -- 2bb
		x"00", -- 2bc
		x"78", -- 2bd
		x"40", -- 2be
		x"70", -- 2bf
		x"40", -- 2c0
		x"78", -- 2c1
		x"00", -- 2c2
		x"0e", -- 2c3
		x"10", -- 2c4
		x"10", -- 2c5
		x"10", -- 2c6
		x"0e", -- 2c7
		x"00", -- 2c8
		x"00", -- 2c9
		x"00", -- 2ca
		x"00", -- 2cb
		x"00", -- 2cc
		x"78", -- 2cd
		x"40", -- 2ce
		x"70", -- 2cf
		x"40", -- 2d0
		x"40", -- 2d1
		x"00", -- 2d2
		x"0e", -- 2d3
		x"10", -- 2d4
		x"0c", -- 2d5
		x"02", -- 2d6
		x"1c", -- 2d7
		x"00", -- 2d8
		x"00", -- 2d9
		x"00", -- 2da
		x"00", -- 2db
		x"00", -- 2dc
		x"38", -- 2dd
		x"40", -- 2de
		x"58", -- 2df
		x"48", -- 2e0
		x"38", -- 2e1
		x"00", -- 2e2
		x"0e", -- 2e3
		x"10", -- 2e4
		x"0c", -- 2e5
		x"02", -- 2e6
		x"1c", -- 2e7
		x"00", -- 2e8
		x"00", -- 2e9
		x"00", -- 2ea
		x"00", -- 2eb
		x"00", -- 2ec
		x"70", -- 2ed
		x"48", -- 2ee
		x"70", -- 2ef
		x"50", -- 2f0
		x"48", -- 2f1
		x"00", -- 2f2
		x"0e", -- 2f3
		x"10", -- 2f4
		x"0c", -- 2f5
		x"02", -- 2f6
		x"1c", -- 2f7
		x"00", -- 2f8
		x"00", -- 2f9
		x"00", -- 2fa
		x"00", -- 2fb
		x"00", -- 2fc
		x"48", -- 2fd
		x"48", -- 2fe
		x"48", -- 2ff
		x"48", -- 300
		x"30", -- 301
		x"00", -- 302
		x"0e", -- 303
		x"10", -- 304
		x"0c", -- 305
		x"02", -- 306
		x"1c", -- 307
		x"00", -- 308
		x"00", -- 309
		x"00", -- 30a
		x"00", -- 30b
		x"00", -- 30c
		x"00", -- 30d
		x"00", -- 30e
		x"00", -- 30f
		x"00", -- 310
		x"00", -- 311
		x"00", -- 312
		x"00", -- 313
		x"00", -- 314
		x"00", -- 315
		x"00", -- 316
		x"00", -- 317
		x"00", -- 318
		x"00", -- 319
		x"00", -- 31a
		x"00", -- 31b
		x"00", -- 31c
		x"00", -- 31d
		x"10", -- 31e
		x"10", -- 31f
		x"10", -- 320
		x"10", -- 321
		x"10", -- 322
		x"10", -- 323
		x"10", -- 324
		x"10", -- 325
		x"00", -- 326
		x"10", -- 327
		x"00", -- 328
		x"00", -- 329
		x"00", -- 32a
		x"00", -- 32b
		x"00", -- 32c
		x"28", -- 32d
		x"28", -- 32e
		x"28", -- 32f
		x"00", -- 330
		x"00", -- 331
		x"00", -- 332
		x"00", -- 333
		x"00", -- 334
		x"00", -- 335
		x"00", -- 336
		x"00", -- 337
		x"00", -- 338
		x"00", -- 339
		x"00", -- 33a
		x"00", -- 33b
		x"00", -- 33c
		x"00", -- 33d
		x"24", -- 33e
		x"24", -- 33f
		x"7e", -- 340
		x"24", -- 341
		x"24", -- 342
		x"24", -- 343
		x"24", -- 344
		x"7e", -- 345
		x"24", -- 346
		x"24", -- 347
		x"00", -- 348
		x"00", -- 349
		x"00", -- 34a
		x"00", -- 34b
		x"00", -- 34c
		x"00", -- 34d
		x"10", -- 34e
		x"38", -- 34f
		x"54", -- 350
		x"50", -- 351
		x"30", -- 352
		x"18", -- 353
		x"14", -- 354
		x"54", -- 355
		x"38", -- 356
		x"10", -- 357
		x"00", -- 358
		x"00", -- 359
		x"00", -- 35a
		x"00", -- 35b
		x"00", -- 35c
		x"00", -- 35d
		x"22", -- 35e
		x"54", -- 35f
		x"24", -- 360
		x"08", -- 361
		x"08", -- 362
		x"10", -- 363
		x"10", -- 364
		x"24", -- 365
		x"2a", -- 366
		x"44", -- 367
		x"00", -- 368
		x"00", -- 369
		x"00", -- 36a
		x"00", -- 36b
		x"00", -- 36c
		x"00", -- 36d
		x"30", -- 36e
		x"48", -- 36f
		x"48", -- 370
		x"50", -- 371
		x"20", -- 372
		x"50", -- 373
		x"8a", -- 374
		x"84", -- 375
		x"8c", -- 376
		x"72", -- 377
		x"00", -- 378
		x"00", -- 379
		x"00", -- 37a
		x"00", -- 37b
		x"00", -- 37c
		x"00", -- 37d
		x"08", -- 37e
		x"10", -- 37f
		x"20", -- 380
		x"00", -- 381
		x"00", -- 382
		x"00", -- 383
		x"00", -- 384
		x"00", -- 385
		x"00", -- 386
		x"00", -- 387
		x"00", -- 388
		x"00", -- 389
		x"00", -- 38a
		x"00", -- 38b
		x"00", -- 38c
		x"00", -- 38d
		x"08", -- 38e
		x"10", -- 38f
		x"10", -- 390
		x"20", -- 391
		x"20", -- 392
		x"20", -- 393
		x"20", -- 394
		x"10", -- 395
		x"10", -- 396
		x"08", -- 397
		x"00", -- 398
		x"00", -- 399
		x"00", -- 39a
		x"00", -- 39b
		x"00", -- 39c
		x"00", -- 39d
		x"20", -- 39e
		x"10", -- 39f
		x"10", -- 3a0
		x"08", -- 3a1
		x"08", -- 3a2
		x"08", -- 3a3
		x"08", -- 3a4
		x"10", -- 3a5
		x"10", -- 3a6
		x"20", -- 3a7
		x"00", -- 3a8
		x"00", -- 3a9
		x"00", -- 3aa
		x"00", -- 3ab
		x"00", -- 3ac
		x"00", -- 3ad
		x"00", -- 3ae
		x"00", -- 3af
		x"10", -- 3b0
		x"54", -- 3b1
		x"38", -- 3b2
		x"38", -- 3b3
		x"54", -- 3b4
		x"10", -- 3b5
		x"00", -- 3b6
		x"00", -- 3b7
		x"00", -- 3b8
		x"00", -- 3b9
		x"00", -- 3ba
		x"00", -- 3bb
		x"00", -- 3bc
		x"00", -- 3bd
		x"00", -- 3be
		x"00", -- 3bf
		x"10", -- 3c0
		x"10", -- 3c1
		x"10", -- 3c2
		x"fe", -- 3c3
		x"10", -- 3c4
		x"10", -- 3c5
		x"10", -- 3c6
		x"00", -- 3c7
		x"00", -- 3c8
		x"00", -- 3c9
		x"00", -- 3ca
		x"00", -- 3cb
		x"00", -- 3cc
		x"00", -- 3cd
		x"00", -- 3ce
		x"00", -- 3cf
		x"00", -- 3d0
		x"00", -- 3d1
		x"00", -- 3d2
		x"00", -- 3d3
		x"00", -- 3d4
		x"00", -- 3d5
		x"30", -- 3d6
		x"30", -- 3d7
		x"10", -- 3d8
		x"20", -- 3d9
		x"00", -- 3da
		x"00", -- 3db
		x"00", -- 3dc
		x"00", -- 3dd
		x"00", -- 3de
		x"00", -- 3df
		x"00", -- 3e0
		x"00", -- 3e1
		x"00", -- 3e2
		x"7e", -- 3e3
		x"00", -- 3e4
		x"00", -- 3e5
		x"00", -- 3e6
		x"00", -- 3e7
		x"00", -- 3e8
		x"00", -- 3e9
		x"00", -- 3ea
		x"00", -- 3eb
		x"00", -- 3ec
		x"00", -- 3ed
		x"00", -- 3ee
		x"00", -- 3ef
		x"00", -- 3f0
		x"00", -- 3f1
		x"00", -- 3f2
		x"00", -- 3f3
		x"00", -- 3f4
		x"00", -- 3f5
		x"30", -- 3f6
		x"30", -- 3f7
		x"00", -- 3f8
		x"00", -- 3f9
		x"00", -- 3fa
		x"00", -- 3fb
		x"00", -- 3fc
		x"00", -- 3fd
		x"04", -- 3fe
		x"04", -- 3ff
		x"08", -- 400
		x"08", -- 401
		x"10", -- 402
		x"10", -- 403
		x"20", -- 404
		x"20", -- 405
		x"40", -- 406
		x"40", -- 407
		x"00", -- 408
		x"00", -- 409
		x"00", -- 40a
		x"00", -- 40b
		x"00", -- 40c
		x"00", -- 40d
		x"3c", -- 40e
		x"42", -- 40f
		x"42", -- 410
		x"46", -- 411
		x"4a", -- 412
		x"52", -- 413
		x"62", -- 414
		x"42", -- 415
		x"42", -- 416
		x"3c", -- 417
		x"00", -- 418
		x"00", -- 419
		x"00", -- 41a
		x"00", -- 41b
		x"00", -- 41c
		x"00", -- 41d
		x"08", -- 41e
		x"18", -- 41f
		x"08", -- 420
		x"08", -- 421
		x"08", -- 422
		x"08", -- 423
		x"08", -- 424
		x"08", -- 425
		x"08", -- 426
		x"1c", -- 427
		x"00", -- 428
		x"00", -- 429
		x"00", -- 42a
		x"00", -- 42b
		x"00", -- 42c
		x"00", -- 42d
		x"3c", -- 42e
		x"42", -- 42f
		x"02", -- 430
		x"02", -- 431
		x"0c", -- 432
		x"10", -- 433
		x"20", -- 434
		x"40", -- 435
		x"40", -- 436
		x"7e", -- 437
		x"00", -- 438
		x"00", -- 439
		x"00", -- 43a
		x"00", -- 43b
		x"00", -- 43c
		x"00", -- 43d
		x"3c", -- 43e
		x"42", -- 43f
		x"02", -- 440
		x"02", -- 441
		x"1c", -- 442
		x"02", -- 443
		x"02", -- 444
		x"02", -- 445
		x"42", -- 446
		x"3c", -- 447
		x"00", -- 448
		x"00", -- 449
		x"00", -- 44a
		x"00", -- 44b
		x"00", -- 44c
		x"00", -- 44d
		x"04", -- 44e
		x"0c", -- 44f
		x"14", -- 450
		x"24", -- 451
		x"44", -- 452
		x"7e", -- 453
		x"04", -- 454
		x"04", -- 455
		x"04", -- 456
		x"04", -- 457
		x"00", -- 458
		x"00", -- 459
		x"00", -- 45a
		x"00", -- 45b
		x"00", -- 45c
		x"00", -- 45d
		x"7c", -- 45e
		x"40", -- 45f
		x"40", -- 460
		x"40", -- 461
		x"7c", -- 462
		x"02", -- 463
		x"02", -- 464
		x"02", -- 465
		x"42", -- 466
		x"3c", -- 467
		x"00", -- 468
		x"00", -- 469
		x"00", -- 46a
		x"00", -- 46b
		x"00", -- 46c
		x"00", -- 46d
		x"3c", -- 46e
		x"42", -- 46f
		x"40", -- 470
		x"40", -- 471
		x"7c", -- 472
		x"42", -- 473
		x"42", -- 474
		x"42", -- 475
		x"42", -- 476
		x"3c", -- 477
		x"00", -- 478
		x"00", -- 479
		x"00", -- 47a
		x"00", -- 47b
		x"00", -- 47c
		x"00", -- 47d
		x"7e", -- 47e
		x"02", -- 47f
		x"02", -- 480
		x"04", -- 481
		x"08", -- 482
		x"08", -- 483
		x"10", -- 484
		x"10", -- 485
		x"20", -- 486
		x"20", -- 487
		x"00", -- 488
		x"00", -- 489
		x"00", -- 48a
		x"00", -- 48b
		x"00", -- 48c
		x"00", -- 48d
		x"3c", -- 48e
		x"42", -- 48f
		x"42", -- 490
		x"42", -- 491
		x"3c", -- 492
		x"42", -- 493
		x"42", -- 494
		x"42", -- 495
		x"42", -- 496
		x"3c", -- 497
		x"00", -- 498
		x"00", -- 499
		x"00", -- 49a
		x"00", -- 49b
		x"00", -- 49c
		x"00", -- 49d
		x"3c", -- 49e
		x"42", -- 49f
		x"42", -- 4a0
		x"42", -- 4a1
		x"3e", -- 4a2
		x"02", -- 4a3
		x"02", -- 4a4
		x"02", -- 4a5
		x"42", -- 4a6
		x"3c", -- 4a7
		x"00", -- 4a8
		x"00", -- 4a9
		x"00", -- 4aa
		x"00", -- 4ab
		x"00", -- 4ac
		x"00", -- 4ad
		x"00", -- 4ae
		x"00", -- 4af
		x"00", -- 4b0
		x"30", -- 4b1
		x"30", -- 4b2
		x"00", -- 4b3
		x"00", -- 4b4
		x"00", -- 4b5
		x"30", -- 4b6
		x"30", -- 4b7
		x"00", -- 4b8
		x"00", -- 4b9
		x"00", -- 4ba
		x"00", -- 4bb
		x"00", -- 4bc
		x"00", -- 4bd
		x"00", -- 4be
		x"00", -- 4bf
		x"00", -- 4c0
		x"30", -- 4c1
		x"30", -- 4c2
		x"00", -- 4c3
		x"00", -- 4c4
		x"00", -- 4c5
		x"30", -- 4c6
		x"30", -- 4c7
		x"10", -- 4c8
		x"20", -- 4c9
		x"00", -- 4ca
		x"00", -- 4cb
		x"00", -- 4cc
		x"00", -- 4cd
		x"00", -- 4ce
		x"08", -- 4cf
		x"10", -- 4d0
		x"20", -- 4d1
		x"40", -- 4d2
		x"20", -- 4d3
		x"10", -- 4d4
		x"08", -- 4d5
		x"00", -- 4d6
		x"00", -- 4d7
		x"00", -- 4d8
		x"00", -- 4d9
		x"00", -- 4da
		x"00", -- 4db
		x"00", -- 4dc
		x"00", -- 4dd
		x"00", -- 4de
		x"00", -- 4df
		x"00", -- 4e0
		x"7e", -- 4e1
		x"00", -- 4e2
		x"00", -- 4e3
		x"7e", -- 4e4
		x"00", -- 4e5
		x"00", -- 4e6
		x"00", -- 4e7
		x"00", -- 4e8
		x"00", -- 4e9
		x"00", -- 4ea
		x"00", -- 4eb
		x"00", -- 4ec
		x"00", -- 4ed
		x"00", -- 4ee
		x"20", -- 4ef
		x"10", -- 4f0
		x"08", -- 4f1
		x"04", -- 4f2
		x"08", -- 4f3
		x"10", -- 4f4
		x"20", -- 4f5
		x"00", -- 4f6
		x"00", -- 4f7
		x"00", -- 4f8
		x"00", -- 4f9
		x"00", -- 4fa
		x"00", -- 4fb
		x"00", -- 4fc
		x"00", -- 4fd
		x"3c", -- 4fe
		x"42", -- 4ff
		x"02", -- 500
		x"02", -- 501
		x"04", -- 502
		x"08", -- 503
		x"10", -- 504
		x"10", -- 505
		x"00", -- 506
		x"10", -- 507
		x"00", -- 508
		x"00", -- 509
		x"00", -- 50a
		x"00", -- 50b
		x"00", -- 50c
		x"00", -- 50d
		x"3c", -- 50e
		x"42", -- 50f
		x"4e", -- 510
		x"52", -- 511
		x"52", -- 512
		x"52", -- 513
		x"4c", -- 514
		x"40", -- 515
		x"42", -- 516
		x"3c", -- 517
		x"00", -- 518
		x"00", -- 519
		x"00", -- 51a
		x"00", -- 51b
		x"00", -- 51c
		x"00", -- 51d
		x"3c", -- 51e
		x"42", -- 51f
		x"42", -- 520
		x"42", -- 521
		x"7e", -- 522
		x"42", -- 523
		x"42", -- 524
		x"42", -- 525
		x"42", -- 526
		x"42", -- 527
		x"00", -- 528
		x"00", -- 529
		x"00", -- 52a
		x"00", -- 52b
		x"00", -- 52c
		x"00", -- 52d
		x"7c", -- 52e
		x"42", -- 52f
		x"42", -- 530
		x"42", -- 531
		x"7c", -- 532
		x"42", -- 533
		x"42", -- 534
		x"42", -- 535
		x"42", -- 536
		x"7c", -- 537
		x"00", -- 538
		x"00", -- 539
		x"00", -- 53a
		x"00", -- 53b
		x"00", -- 53c
		x"00", -- 53d
		x"3c", -- 53e
		x"42", -- 53f
		x"40", -- 540
		x"40", -- 541
		x"40", -- 542
		x"40", -- 543
		x"40", -- 544
		x"40", -- 545
		x"42", -- 546
		x"3c", -- 547
		x"00", -- 548
		x"00", -- 549
		x"00", -- 54a
		x"00", -- 54b
		x"00", -- 54c
		x"00", -- 54d
		x"7c", -- 54e
		x"42", -- 54f
		x"42", -- 550
		x"42", -- 551
		x"42", -- 552
		x"42", -- 553
		x"42", -- 554
		x"42", -- 555
		x"42", -- 556
		x"7c", -- 557
		x"00", -- 558
		x"00", -- 559
		x"00", -- 55a
		x"00", -- 55b
		x"00", -- 55c
		x"00", -- 55d
		x"7e", -- 55e
		x"40", -- 55f
		x"40", -- 560
		x"40", -- 561
		x"7c", -- 562
		x"40", -- 563
		x"40", -- 564
		x"40", -- 565
		x"40", -- 566
		x"7e", -- 567
		x"00", -- 568
		x"00", -- 569
		x"00", -- 56a
		x"00", -- 56b
		x"00", -- 56c
		x"00", -- 56d
		x"7e", -- 56e
		x"40", -- 56f
		x"40", -- 570
		x"40", -- 571
		x"78", -- 572
		x"40", -- 573
		x"40", -- 574
		x"40", -- 575
		x"40", -- 576
		x"40", -- 577
		x"00", -- 578
		x"00", -- 579
		x"00", -- 57a
		x"00", -- 57b
		x"00", -- 57c
		x"00", -- 57d
		x"3c", -- 57e
		x"42", -- 57f
		x"40", -- 580
		x"40", -- 581
		x"40", -- 582
		x"4e", -- 583
		x"42", -- 584
		x"42", -- 585
		x"42", -- 586
		x"3c", -- 587
		x"00", -- 588
		x"00", -- 589
		x"00", -- 58a
		x"00", -- 58b
		x"00", -- 58c
		x"00", -- 58d
		x"42", -- 58e
		x"42", -- 58f
		x"42", -- 590
		x"42", -- 591
		x"7e", -- 592
		x"42", -- 593
		x"42", -- 594
		x"42", -- 595
		x"42", -- 596
		x"42", -- 597
		x"00", -- 598
		x"00", -- 599
		x"00", -- 59a
		x"00", -- 59b
		x"00", -- 59c
		x"00", -- 59d
		x"38", -- 59e
		x"10", -- 59f
		x"10", -- 5a0
		x"10", -- 5a1
		x"10", -- 5a2
		x"10", -- 5a3
		x"10", -- 5a4
		x"10", -- 5a5
		x"10", -- 5a6
		x"38", -- 5a7
		x"00", -- 5a8
		x"00", -- 5a9
		x"00", -- 5aa
		x"00", -- 5ab
		x"00", -- 5ac
		x"00", -- 5ad
		x"0e", -- 5ae
		x"04", -- 5af
		x"04", -- 5b0
		x"04", -- 5b1
		x"04", -- 5b2
		x"04", -- 5b3
		x"04", -- 5b4
		x"04", -- 5b5
		x"44", -- 5b6
		x"38", -- 5b7
		x"00", -- 5b8
		x"00", -- 5b9
		x"00", -- 5ba
		x"00", -- 5bb
		x"00", -- 5bc
		x"00", -- 5bd
		x"42", -- 5be
		x"44", -- 5bf
		x"48", -- 5c0
		x"50", -- 5c1
		x"60", -- 5c2
		x"50", -- 5c3
		x"48", -- 5c4
		x"44", -- 5c5
		x"42", -- 5c6
		x"42", -- 5c7
		x"00", -- 5c8
		x"00", -- 5c9
		x"00", -- 5ca
		x"00", -- 5cb
		x"00", -- 5cc
		x"00", -- 5cd
		x"40", -- 5ce
		x"40", -- 5cf
		x"40", -- 5d0
		x"40", -- 5d1
		x"40", -- 5d2
		x"40", -- 5d3
		x"40", -- 5d4
		x"40", -- 5d5
		x"40", -- 5d6
		x"7e", -- 5d7
		x"00", -- 5d8
		x"00", -- 5d9
		x"00", -- 5da
		x"00", -- 5db
		x"00", -- 5dc
		x"00", -- 5dd
		x"82", -- 5de
		x"82", -- 5df
		x"c6", -- 5e0
		x"aa", -- 5e1
		x"92", -- 5e2
		x"82", -- 5e3
		x"82", -- 5e4
		x"82", -- 5e5
		x"82", -- 5e6
		x"82", -- 5e7
		x"00", -- 5e8
		x"00", -- 5e9
		x"00", -- 5ea
		x"00", -- 5eb
		x"00", -- 5ec
		x"00", -- 5ed
		x"42", -- 5ee
		x"62", -- 5ef
		x"62", -- 5f0
		x"52", -- 5f1
		x"52", -- 5f2
		x"4a", -- 5f3
		x"4a", -- 5f4
		x"46", -- 5f5
		x"46", -- 5f6
		x"42", -- 5f7
		x"00", -- 5f8
		x"00", -- 5f9
		x"00", -- 5fa
		x"00", -- 5fb
		x"00", -- 5fc
		x"00", -- 5fd
		x"3c", -- 5fe
		x"42", -- 5ff
		x"42", -- 600
		x"42", -- 601
		x"42", -- 602
		x"42", -- 603
		x"42", -- 604
		x"42", -- 605
		x"42", -- 606
		x"3c", -- 607
		x"00", -- 608
		x"00", -- 609
		x"00", -- 60a
		x"00", -- 60b
		x"00", -- 60c
		x"00", -- 60d
		x"7c", -- 60e
		x"42", -- 60f
		x"42", -- 610
		x"42", -- 611
		x"7c", -- 612
		x"40", -- 613
		x"40", -- 614
		x"40", -- 615
		x"40", -- 616
		x"40", -- 617
		x"00", -- 618
		x"00", -- 619
		x"00", -- 61a
		x"00", -- 61b
		x"00", -- 61c
		x"00", -- 61d
		x"3c", -- 61e
		x"42", -- 61f
		x"42", -- 620
		x"42", -- 621
		x"42", -- 622
		x"42", -- 623
		x"42", -- 624
		x"42", -- 625
		x"4a", -- 626
		x"3c", -- 627
		x"04", -- 628
		x"02", -- 629
		x"00", -- 62a
		x"00", -- 62b
		x"00", -- 62c
		x"00", -- 62d
		x"7c", -- 62e
		x"42", -- 62f
		x"42", -- 630
		x"42", -- 631
		x"7c", -- 632
		x"48", -- 633
		x"44", -- 634
		x"42", -- 635
		x"42", -- 636
		x"42", -- 637
		x"00", -- 638
		x"00", -- 639
		x"00", -- 63a
		x"00", -- 63b
		x"00", -- 63c
		x"00", -- 63d
		x"3c", -- 63e
		x"42", -- 63f
		x"40", -- 640
		x"40", -- 641
		x"3c", -- 642
		x"02", -- 643
		x"02", -- 644
		x"02", -- 645
		x"42", -- 646
		x"3c", -- 647
		x"00", -- 648
		x"00", -- 649
		x"00", -- 64a
		x"00", -- 64b
		x"00", -- 64c
		x"00", -- 64d
		x"fe", -- 64e
		x"10", -- 64f
		x"10", -- 650
		x"10", -- 651
		x"10", -- 652
		x"10", -- 653
		x"10", -- 654
		x"10", -- 655
		x"10", -- 656
		x"10", -- 657
		x"00", -- 658
		x"00", -- 659
		x"00", -- 65a
		x"00", -- 65b
		x"00", -- 65c
		x"00", -- 65d
		x"42", -- 65e
		x"42", -- 65f
		x"42", -- 660
		x"42", -- 661
		x"42", -- 662
		x"42", -- 663
		x"42", -- 664
		x"42", -- 665
		x"42", -- 666
		x"3c", -- 667
		x"00", -- 668
		x"00", -- 669
		x"00", -- 66a
		x"00", -- 66b
		x"00", -- 66c
		x"00", -- 66d
		x"82", -- 66e
		x"82", -- 66f
		x"44", -- 670
		x"44", -- 671
		x"44", -- 672
		x"28", -- 673
		x"28", -- 674
		x"28", -- 675
		x"10", -- 676
		x"10", -- 677
		x"00", -- 678
		x"00", -- 679
		x"00", -- 67a
		x"00", -- 67b
		x"00", -- 67c
		x"00", -- 67d
		x"82", -- 67e
		x"82", -- 67f
		x"82", -- 680
		x"82", -- 681
		x"82", -- 682
		x"92", -- 683
		x"aa", -- 684
		x"c6", -- 685
		x"82", -- 686
		x"82", -- 687
		x"00", -- 688
		x"00", -- 689
		x"00", -- 68a
		x"00", -- 68b
		x"00", -- 68c
		x"00", -- 68d
		x"42", -- 68e
		x"42", -- 68f
		x"42", -- 690
		x"24", -- 691
		x"18", -- 692
		x"18", -- 693
		x"24", -- 694
		x"42", -- 695
		x"42", -- 696
		x"42", -- 697
		x"00", -- 698
		x"00", -- 699
		x"00", -- 69a
		x"00", -- 69b
		x"00", -- 69c
		x"00", -- 69d
		x"82", -- 69e
		x"82", -- 69f
		x"44", -- 6a0
		x"44", -- 6a1
		x"28", -- 6a2
		x"10", -- 6a3
		x"10", -- 6a4
		x"10", -- 6a5
		x"10", -- 6a6
		x"10", -- 6a7
		x"00", -- 6a8
		x"00", -- 6a9
		x"00", -- 6aa
		x"00", -- 6ab
		x"00", -- 6ac
		x"00", -- 6ad
		x"7e", -- 6ae
		x"02", -- 6af
		x"02", -- 6b0
		x"04", -- 6b1
		x"08", -- 6b2
		x"10", -- 6b3
		x"20", -- 6b4
		x"40", -- 6b5
		x"40", -- 6b6
		x"7e", -- 6b7
		x"00", -- 6b8
		x"00", -- 6b9
		x"00", -- 6ba
		x"00", -- 6bb
		x"00", -- 6bc
		x"00", -- 6bd
		x"3c", -- 6be
		x"20", -- 6bf
		x"20", -- 6c0
		x"20", -- 6c1
		x"20", -- 6c2
		x"20", -- 6c3
		x"20", -- 6c4
		x"20", -- 6c5
		x"20", -- 6c6
		x"3c", -- 6c7
		x"00", -- 6c8
		x"00", -- 6c9
		x"00", -- 6ca
		x"00", -- 6cb
		x"00", -- 6cc
		x"00", -- 6cd
		x"40", -- 6ce
		x"40", -- 6cf
		x"20", -- 6d0
		x"20", -- 6d1
		x"10", -- 6d2
		x"10", -- 6d3
		x"08", -- 6d4
		x"08", -- 6d5
		x"04", -- 6d6
		x"04", -- 6d7
		x"00", -- 6d8
		x"00", -- 6d9
		x"00", -- 6da
		x"00", -- 6db
		x"00", -- 6dc
		x"00", -- 6dd
		x"3c", -- 6de
		x"04", -- 6df
		x"04", -- 6e0
		x"04", -- 6e1
		x"04", -- 6e2
		x"04", -- 6e3
		x"04", -- 6e4
		x"04", -- 6e5
		x"04", -- 6e6
		x"3c", -- 6e7
		x"00", -- 6e8
		x"00", -- 6e9
		x"00", -- 6ea
		x"00", -- 6eb
		x"00", -- 6ec
		x"00", -- 6ed
		x"10", -- 6ee
		x"28", -- 6ef
		x"44", -- 6f0
		x"00", -- 6f1
		x"00", -- 6f2
		x"00", -- 6f3
		x"00", -- 6f4
		x"00", -- 6f5
		x"00", -- 6f6
		x"00", -- 6f7
		x"00", -- 6f8
		x"00", -- 6f9
		x"00", -- 6fa
		x"00", -- 6fb
		x"00", -- 6fc
		x"00", -- 6fd
		x"00", -- 6fe
		x"00", -- 6ff
		x"00", -- 700
		x"00", -- 701
		x"00", -- 702
		x"00", -- 703
		x"00", -- 704
		x"00", -- 705
		x"00", -- 706
		x"00", -- 707
		x"00", -- 708
		x"ff", -- 709
		x"00", -- 70a
		x"00", -- 70b
		x"00", -- 70c
		x"20", -- 70d
		x"10", -- 70e
		x"08", -- 70f
		x"04", -- 710
		x"00", -- 711
		x"00", -- 712
		x"00", -- 713
		x"00", -- 714
		x"00", -- 715
		x"00", -- 716
		x"00", -- 717
		x"00", -- 718
		x"00", -- 719
		x"00", -- 71a
		x"00", -- 71b
		x"00", -- 71c
		x"00", -- 71d
		x"00", -- 71e
		x"00", -- 71f
		x"00", -- 720
		x"00", -- 721
		x"3c", -- 722
		x"02", -- 723
		x"3e", -- 724
		x"42", -- 725
		x"42", -- 726
		x"3e", -- 727
		x"00", -- 728
		x"00", -- 729
		x"00", -- 72a
		x"00", -- 72b
		x"00", -- 72c
		x"00", -- 72d
		x"40", -- 72e
		x"40", -- 72f
		x"40", -- 730
		x"40", -- 731
		x"7c", -- 732
		x"42", -- 733
		x"42", -- 734
		x"42", -- 735
		x"42", -- 736
		x"7c", -- 737
		x"00", -- 738
		x"00", -- 739
		x"00", -- 73a
		x"00", -- 73b
		x"00", -- 73c
		x"00", -- 73d
		x"00", -- 73e
		x"00", -- 73f
		x"00", -- 740
		x"00", -- 741
		x"3c", -- 742
		x"42", -- 743
		x"40", -- 744
		x"40", -- 745
		x"42", -- 746
		x"3c", -- 747
		x"00", -- 748
		x"00", -- 749
		x"00", -- 74a
		x"00", -- 74b
		x"00", -- 74c
		x"00", -- 74d
		x"02", -- 74e
		x"02", -- 74f
		x"02", -- 750
		x"02", -- 751
		x"3e", -- 752
		x"42", -- 753
		x"42", -- 754
		x"42", -- 755
		x"42", -- 756
		x"3e", -- 757
		x"00", -- 758
		x"00", -- 759
		x"00", -- 75a
		x"00", -- 75b
		x"00", -- 75c
		x"00", -- 75d
		x"00", -- 75e
		x"00", -- 75f
		x"00", -- 760
		x"00", -- 761
		x"3c", -- 762
		x"42", -- 763
		x"7e", -- 764
		x"40", -- 765
		x"42", -- 766
		x"3c", -- 767
		x"00", -- 768
		x"00", -- 769
		x"00", -- 76a
		x"00", -- 76b
		x"00", -- 76c
		x"00", -- 76d
		x"18", -- 76e
		x"24", -- 76f
		x"20", -- 770
		x"20", -- 771
		x"20", -- 772
		x"78", -- 773
		x"20", -- 774
		x"20", -- 775
		x"20", -- 776
		x"20", -- 777
		x"00", -- 778
		x"00", -- 779
		x"00", -- 77a
		x"00", -- 77b
		x"00", -- 77c
		x"00", -- 77d
		x"00", -- 77e
		x"00", -- 77f
		x"00", -- 780
		x"00", -- 781
		x"3e", -- 782
		x"42", -- 783
		x"42", -- 784
		x"42", -- 785
		x"42", -- 786
		x"3e", -- 787
		x"02", -- 788
		x"02", -- 789
		x"3c", -- 78a
		x"00", -- 78b
		x"00", -- 78c
		x"00", -- 78d
		x"40", -- 78e
		x"40", -- 78f
		x"40", -- 790
		x"40", -- 791
		x"7c", -- 792
		x"42", -- 793
		x"42", -- 794
		x"42", -- 795
		x"42", -- 796
		x"42", -- 797
		x"00", -- 798
		x"00", -- 799
		x"00", -- 79a
		x"00", -- 79b
		x"00", -- 79c
		x"00", -- 79d
		x"00", -- 79e
		x"00", -- 79f
		x"10", -- 7a0
		x"00", -- 7a1
		x"30", -- 7a2
		x"10", -- 7a3
		x"10", -- 7a4
		x"10", -- 7a5
		x"10", -- 7a6
		x"38", -- 7a7
		x"00", -- 7a8
		x"00", -- 7a9
		x"00", -- 7aa
		x"00", -- 7ab
		x"00", -- 7ac
		x"00", -- 7ad
		x"00", -- 7ae
		x"00", -- 7af
		x"04", -- 7b0
		x"00", -- 7b1
		x"0c", -- 7b2
		x"04", -- 7b3
		x"04", -- 7b4
		x"04", -- 7b5
		x"04", -- 7b6
		x"04", -- 7b7
		x"04", -- 7b8
		x"04", -- 7b9
		x"18", -- 7ba
		x"00", -- 7bb
		x"00", -- 7bc
		x"00", -- 7bd
		x"40", -- 7be
		x"40", -- 7bf
		x"40", -- 7c0
		x"40", -- 7c1
		x"44", -- 7c2
		x"48", -- 7c3
		x"50", -- 7c4
		x"68", -- 7c5
		x"44", -- 7c6
		x"44", -- 7c7
		x"00", -- 7c8
		x"00", -- 7c9
		x"00", -- 7ca
		x"00", -- 7cb
		x"00", -- 7cc
		x"00", -- 7cd
		x"18", -- 7ce
		x"08", -- 7cf
		x"08", -- 7d0
		x"08", -- 7d1
		x"08", -- 7d2
		x"08", -- 7d3
		x"08", -- 7d4
		x"08", -- 7d5
		x"08", -- 7d6
		x"1c", -- 7d7
		x"00", -- 7d8
		x"00", -- 7d9
		x"00", -- 7da
		x"00", -- 7db
		x"00", -- 7dc
		x"00", -- 7dd
		x"00", -- 7de
		x"00", -- 7df
		x"00", -- 7e0
		x"00", -- 7e1
		x"ec", -- 7e2
		x"92", -- 7e3
		x"92", -- 7e4
		x"92", -- 7e5
		x"92", -- 7e6
		x"92", -- 7e7
		x"00", -- 7e8
		x"00", -- 7e9
		x"00", -- 7ea
		x"00", -- 7eb
		x"00", -- 7ec
		x"00", -- 7ed
		x"00", -- 7ee
		x"00", -- 7ef
		x"00", -- 7f0
		x"00", -- 7f1
		x"5c", -- 7f2
		x"62", -- 7f3
		x"42", -- 7f4
		x"42", -- 7f5
		x"42", -- 7f6
		x"42", -- 7f7
		x"00", -- 7f8
		x"00", -- 7f9
		x"00", -- 7fa
		x"00", -- 7fb
		x"00", -- 7fc
		x"00", -- 7fd
		x"00", -- 7fe
		x"00", -- 7ff
		x"00", -- 800
		x"00", -- 801
		x"3c", -- 802
		x"42", -- 803
		x"42", -- 804
		x"42", -- 805
		x"42", -- 806
		x"3c", -- 807
		x"00", -- 808
		x"00", -- 809
		x"00", -- 80a
		x"00", -- 80b
		x"00", -- 80c
		x"00", -- 80d
		x"00", -- 80e
		x"00", -- 80f
		x"00", -- 810
		x"00", -- 811
		x"5c", -- 812
		x"62", -- 813
		x"42", -- 814
		x"42", -- 815
		x"42", -- 816
		x"7c", -- 817
		x"40", -- 818
		x"40", -- 819
		x"40", -- 81a
		x"00", -- 81b
		x"00", -- 81c
		x"00", -- 81d
		x"00", -- 81e
		x"00", -- 81f
		x"00", -- 820
		x"00", -- 821
		x"3a", -- 822
		x"46", -- 823
		x"42", -- 824
		x"42", -- 825
		x"42", -- 826
		x"3e", -- 827
		x"02", -- 828
		x"02", -- 829
		x"02", -- 82a
		x"00", -- 82b
		x"00", -- 82c
		x"00", -- 82d
		x"00", -- 82e
		x"00", -- 82f
		x"00", -- 830
		x"00", -- 831
		x"6c", -- 832
		x"32", -- 833
		x"20", -- 834
		x"20", -- 835
		x"20", -- 836
		x"20", -- 837
		x"00", -- 838
		x"00", -- 839
		x"00", -- 83a
		x"00", -- 83b
		x"00", -- 83c
		x"00", -- 83d
		x"00", -- 83e
		x"00", -- 83f
		x"00", -- 840
		x"00", -- 841
		x"3c", -- 842
		x"40", -- 843
		x"3c", -- 844
		x"02", -- 845
		x"42", -- 846
		x"3c", -- 847
		x"00", -- 848
		x"00", -- 849
		x"00", -- 84a
		x"00", -- 84b
		x"00", -- 84c
		x"00", -- 84d
		x"00", -- 84e
		x"00", -- 84f
		x"00", -- 850
		x"10", -- 851
		x"7c", -- 852
		x"10", -- 853
		x"10", -- 854
		x"10", -- 855
		x"10", -- 856
		x"0c", -- 857
		x"00", -- 858
		x"00", -- 859
		x"00", -- 85a
		x"00", -- 85b
		x"00", -- 85c
		x"00", -- 85d
		x"00", -- 85e
		x"00", -- 85f
		x"00", -- 860
		x"00", -- 861
		x"42", -- 862
		x"42", -- 863
		x"42", -- 864
		x"42", -- 865
		x"42", -- 866
		x"3e", -- 867
		x"00", -- 868
		x"00", -- 869
		x"00", -- 86a
		x"00", -- 86b
		x"00", -- 86c
		x"00", -- 86d
		x"00", -- 86e
		x"00", -- 86f
		x"00", -- 870
		x"00", -- 871
		x"82", -- 872
		x"44", -- 873
		x"44", -- 874
		x"28", -- 875
		x"28", -- 876
		x"10", -- 877
		x"00", -- 878
		x"00", -- 879
		x"00", -- 87a
		x"00", -- 87b
		x"00", -- 87c
		x"00", -- 87d
		x"00", -- 87e
		x"00", -- 87f
		x"00", -- 880
		x"00", -- 881
		x"92", -- 882
		x"92", -- 883
		x"92", -- 884
		x"92", -- 885
		x"92", -- 886
		x"6c", -- 887
		x"00", -- 888
		x"00", -- 889
		x"00", -- 88a
		x"00", -- 88b
		x"00", -- 88c
		x"00", -- 88d
		x"00", -- 88e
		x"00", -- 88f
		x"00", -- 890
		x"00", -- 891
		x"42", -- 892
		x"24", -- 893
		x"18", -- 894
		x"18", -- 895
		x"24", -- 896
		x"42", -- 897
		x"00", -- 898
		x"00", -- 899
		x"00", -- 89a
		x"00", -- 89b
		x"00", -- 89c
		x"00", -- 89d
		x"00", -- 89e
		x"00", -- 89f
		x"00", -- 8a0
		x"00", -- 8a1
		x"42", -- 8a2
		x"42", -- 8a3
		x"42", -- 8a4
		x"42", -- 8a5
		x"42", -- 8a6
		x"3e", -- 8a7
		x"02", -- 8a8
		x"02", -- 8a9
		x"3c", -- 8aa
		x"00", -- 8ab
		x"00", -- 8ac
		x"00", -- 8ad
		x"00", -- 8ae
		x"00", -- 8af
		x"00", -- 8b0
		x"00", -- 8b1
		x"7e", -- 8b2
		x"04", -- 8b3
		x"08", -- 8b4
		x"10", -- 8b5
		x"20", -- 8b6
		x"7e", -- 8b7
		x"00", -- 8b8
		x"00", -- 8b9
		x"00", -- 8ba
		x"00", -- 8bb
		x"00", -- 8bc
		x"00", -- 8bd
		x"0c", -- 8be
		x"10", -- 8bf
		x"10", -- 8c0
		x"10", -- 8c1
		x"10", -- 8c2
		x"20", -- 8c3
		x"10", -- 8c4
		x"10", -- 8c5
		x"10", -- 8c6
		x"0c", -- 8c7
		x"00", -- 8c8
		x"00", -- 8c9
		x"00", -- 8ca
		x"00", -- 8cb
		x"10", -- 8cc
		x"10", -- 8cd
		x"10", -- 8ce
		x"10", -- 8cf
		x"10", -- 8d0
		x"10", -- 8d1
		x"10", -- 8d2
		x"10", -- 8d3
		x"10", -- 8d4
		x"10", -- 8d5
		x"10", -- 8d6
		x"10", -- 8d7
		x"10", -- 8d8
		x"10", -- 8d9
		x"10", -- 8da
		x"10", -- 8db
		x"00", -- 8dc
		x"00", -- 8dd
		x"30", -- 8de
		x"08", -- 8df
		x"08", -- 8e0
		x"08", -- 8e1
		x"08", -- 8e2
		x"04", -- 8e3
		x"08", -- 8e4
		x"08", -- 8e5
		x"08", -- 8e6
		x"30", -- 8e7
		x"00", -- 8e8
		x"00", -- 8e9
		x"00", -- 8ea
		x"00", -- 8eb
		x"00", -- 8ec
		x"00", -- 8ed
		x"00", -- 8ee
		x"00", -- 8ef
		x"00", -- 8f0
		x"00", -- 8f1
		x"32", -- 8f2
		x"4c", -- 8f3
		x"00", -- 8f4
		x"00", -- 8f5
		x"00", -- 8f6
		x"00", -- 8f7
		x"00", -- 8f8
		x"00", -- 8f9
		x"00", -- 8fa
		x"00", -- 8fb
		x"00", -- 8fc
		x"00", -- 8fd
		x"2a", -- 8fe
		x"54", -- 8ff
		x"2a", -- 900
		x"54", -- 901
		x"2a", -- 902
		x"54", -- 903
		x"2a", -- 904
		x"54", -- 905
		x"2a", -- 906
		x"54", -- 907
		x"00", -- 908
		x"00", -- 909
		x"00", -- 90a
		x"00", -- 90b
		x"00", -- 90c
		x"38", -- 90d
		x"40", -- 90e
		x"40", -- 90f
		x"40", -- 910
		x"38", -- 911
		x"00", -- 912
		x"10", -- 913
		x"10", -- 914
		x"10", -- 915
		x"10", -- 916
		x"1e", -- 917
		x"00", -- 918
		x"00", -- 919
		x"00", -- 91a
		x"00", -- 91b
		x"00", -- 91c
		x"70", -- 91d
		x"20", -- 91e
		x"20", -- 91f
		x"20", -- 920
		x"70", -- 921
		x"00", -- 922
		x"22", -- 923
		x"22", -- 924
		x"14", -- 925
		x"14", -- 926
		x"08", -- 927
		x"00", -- 928
		x"00", -- 929
		x"00", -- 92a
		x"00", -- 92b
		x"00", -- 92c
		x"70", -- 92d
		x"48", -- 92e
		x"70", -- 92f
		x"48", -- 930
		x"70", -- 931
		x"00", -- 932
		x"0c", -- 933
		x"10", -- 934
		x"16", -- 935
		x"12", -- 936
		x"0c", -- 937
		x"00", -- 938
		x"00", -- 939
		x"00", -- 93a
		x"00", -- 93b
		x"00", -- 93c
		x"70", -- 93d
		x"20", -- 93e
		x"20", -- 93f
		x"20", -- 940
		x"70", -- 941
		x"00", -- 942
		x"1c", -- 943
		x"12", -- 944
		x"1c", -- 945
		x"12", -- 946
		x"1c", -- 947
		x"00", -- 948
		x"00", -- 949
		x"00", -- 94a
		x"00", -- 94b
		x"00", -- 94c
		x"48", -- 94d
		x"48", -- 94e
		x"48", -- 94f
		x"48", -- 950
		x"30", -- 951
		x"00", -- 952
		x"10", -- 953
		x"10", -- 954
		x"10", -- 955
		x"10", -- 956
		x"1e", -- 957
		x"00", -- 958
		x"ff", -- 959
		x"00", -- 95a
		x"00", -- 95b
		x"00", -- 95c
		x"70", -- 95d
		x"20", -- 95e
		x"20", -- 95f
		x"20", -- 960
		x"70", -- 961
		x"00", -- 962
		x"22", -- 963
		x"22", -- 964
		x"14", -- 965
		x"14", -- 966
		x"08", -- 967
		x"00", -- 968
		x"ff", -- 969
		x"00", -- 96a
		x"00", -- 96b
		x"00", -- 96c
		x"70", -- 96d
		x"48", -- 96e
		x"70", -- 96f
		x"48", -- 970
		x"70", -- 971
		x"00", -- 972
		x"0c", -- 973
		x"10", -- 974
		x"16", -- 975
		x"12", -- 976
		x"0c", -- 977
		x"00", -- 978
		x"ff", -- 979
		x"00", -- 97a
		x"00", -- 97b
		x"00", -- 97c
		x"70", -- 97d
		x"20", -- 97e
		x"20", -- 97f
		x"20", -- 980
		x"70", -- 981
		x"00", -- 982
		x"1c", -- 983
		x"12", -- 984
		x"1c", -- 985
		x"12", -- 986
		x"1c", -- 987
		x"00", -- 988
		x"ff", -- 989
		x"00", -- 98a
		x"00", -- 98b
		x"00", -- 98c
		x"a8", -- 98d
		x"a8", -- 98e
		x"a8", -- 98f
		x"a8", -- 990
		x"50", -- 991
		x"00", -- 992
		x"12", -- 993
		x"12", -- 994
		x"1e", -- 995
		x"12", -- 996
		x"12", -- 997
		x"00", -- 998
		x"00", -- 999
		x"00", -- 99a
		x"00", -- 99b
		x"00", -- 99c
		x"70", -- 99d
		x"48", -- 99e
		x"70", -- 99f
		x"50", -- 9a0
		x"48", -- 9a1
		x"00", -- 9a2
		x"1c", -- 9a3
		x"12", -- 9a4
		x"12", -- 9a5
		x"12", -- 9a6
		x"1c", -- 9a7
		x"00", -- 9a8
		x"00", -- 9a9
		x"00", -- 9aa
		x"00", -- 9ab
		x"00", -- 9ac
		x"44", -- 9ad
		x"28", -- 9ae
		x"10", -- 9af
		x"10", -- 9b0
		x"10", -- 9b1
		x"00", -- 9b2
		x"1e", -- 9b3
		x"10", -- 9b4
		x"1c", -- 9b5
		x"10", -- 9b6
		x"1e", -- 9b7
		x"00", -- 9b8
		x"00", -- 9b9
		x"00", -- 9ba
		x"00", -- 9bb
		x"00", -- 9bc
		x"30", -- 9bd
		x"40", -- 9be
		x"58", -- 9bf
		x"48", -- 9c0
		x"30", -- 9c1
		x"00", -- 9c2
		x"1c", -- 9c3
		x"12", -- 9c4
		x"1c", -- 9c5
		x"14", -- 9c6
		x"12", -- 9c7
		x"00", -- 9c8
		x"00", -- 9c9
		x"00", -- 9ca
		x"00", -- 9cb
		x"00", -- 9cc
		x"38", -- 9cd
		x"40", -- 9ce
		x"40", -- 9cf
		x"40", -- 9d0
		x"38", -- 9d1
		x"00", -- 9d2
		x"22", -- 9d3
		x"14", -- 9d4
		x"08", -- 9d5
		x"08", -- 9d6
		x"08", -- 9d7
		x"00", -- 9d8
		x"00", -- 9d9
		x"00", -- 9da
		x"00", -- 9db
		x"00", -- 9dc
		x"70", -- 9dd
		x"48", -- 9de
		x"70", -- 9df
		x"48", -- 9e0
		x"70", -- 9e1
		x"00", -- 9e2
		x"12", -- 9e3
		x"12", -- 9e4
		x"12", -- 9e5
		x"12", -- 9e6
		x"0c", -- 9e7
		x"00", -- 9e8
		x"00", -- 9e9
		x"00", -- 9ea
		x"00", -- 9eb
		x"00", -- 9ec
		x"88", -- 9ed
		x"d8", -- 9ee
		x"a8", -- 9ef
		x"88", -- 9f0
		x"88", -- 9f1
		x"00", -- 9f2
		x"0c", -- 9f3
		x"10", -- 9f4
		x"16", -- 9f5
		x"12", -- 9f6
		x"0c", -- 9f7
		x"00", -- 9f8
		x"00", -- 9f9
		x"00", -- 9fa
		x"00", -- 9fb
		x"00", -- 9fc
		x"70", -- 9fd
		x"48", -- 9fe
		x"70", -- 9ff
		x"48", -- a00
		x"70", -- a01
		x"00", -- a02
		x"12", -- a03
		x"14", -- a04
		x"18", -- a05
		x"14", -- a06
		x"12", -- a07
		x"00", -- a08
		x"00", -- a09
		x"00", -- a0a
		x"00", -- a0b
		x"00", -- a0c
		x"30", -- a0d
		x"48", -- a0e
		x"38", -- a0f
		x"08", -- a10
		x"30", -- a11
		x"00", -- a12
		x"0c", -- a13
		x"12", -- a14
		x"12", -- a15
		x"12", -- a16
		x"0c", -- a17
		x"00", -- a18
		x"00", -- a19
		x"00", -- a1a
		x"00", -- a1b
		x"00", -- a1c
		x"30", -- a1d
		x"48", -- a1e
		x"38", -- a1f
		x"08", -- a20
		x"30", -- a21
		x"00", -- a22
		x"04", -- a23
		x"0c", -- a24
		x"04", -- a25
		x"04", -- a26
		x"0e", -- a27
		x"00", -- a28
		x"00", -- a29
		x"00", -- a2a
		x"00", -- a2b
		x"00", -- a2c
		x"30", -- a2d
		x"48", -- a2e
		x"38", -- a2f
		x"08", -- a30
		x"30", -- a31
		x"00", -- a32
		x"0c", -- a33
		x"12", -- a34
		x"04", -- a35
		x"08", -- a36
		x"1e", -- a37
		x"00", -- a38
		x"00", -- a39
		x"00", -- a3a
		x"00", -- a3b
		x"00", -- a3c
		x"30", -- a3d
		x"48", -- a3e
		x"38", -- a3f
		x"08", -- a40
		x"30", -- a41
		x"00", -- a42
		x"1c", -- a43
		x"02", -- a44
		x"1c", -- a45
		x"02", -- a46
		x"1c", -- a47
		x"00", -- a48
		x"00", -- a49
		x"00", -- a4a
		x"00", -- a4b
		x"00", -- a4c
		x"30", -- a4d
		x"48", -- a4e
		x"38", -- a4f
		x"08", -- a50
		x"30", -- a51
		x"00", -- a52
		x"14", -- a53
		x"14", -- a54
		x"1e", -- a55
		x"04", -- a56
		x"04", -- a57
		x"00", -- a58
		x"00", -- a59
		x"00", -- a5a
		x"00", -- a5b
		x"00", -- a5c
		x"30", -- a5d
		x"48", -- a5e
		x"38", -- a5f
		x"08", -- a60
		x"30", -- a61
		x"00", -- a62
		x"1e", -- a63
		x"10", -- a64
		x"1c", -- a65
		x"02", -- a66
		x"1c", -- a67
		x"00", -- a68
		x"00", -- a69
		x"00", -- a6a
		x"00", -- a6b
		x"00", -- a6c
		x"30", -- a6d
		x"48", -- a6e
		x"38", -- a6f
		x"08", -- a70
		x"30", -- a71
		x"00", -- a72
		x"0c", -- a73
		x"10", -- a74
		x"1c", -- a75
		x"12", -- a76
		x"0c", -- a77
		x"00", -- a78
		x"00", -- a79
		x"00", -- a7a
		x"00", -- a7b
		x"00", -- a7c
		x"30", -- a7d
		x"48", -- a7e
		x"38", -- a7f
		x"08", -- a80
		x"30", -- a81
		x"00", -- a82
		x"1e", -- a83
		x"02", -- a84
		x"04", -- a85
		x"08", -- a86
		x"10", -- a87
		x"00", -- a88
		x"00", -- a89
		x"00", -- a8a
		x"00", -- a8b
		x"00", -- a8c
		x"30", -- a8d
		x"48", -- a8e
		x"38", -- a8f
		x"08", -- a90
		x"30", -- a91
		x"00", -- a92
		x"0c", -- a93
		x"12", -- a94
		x"0c", -- a95
		x"12", -- a96
		x"0c", -- a97
		x"00", -- a98
		x"00", -- a99
		x"00", -- a9a
		x"00", -- a9b
		x"00", -- a9c
		x"30", -- a9d
		x"48", -- a9e
		x"38", -- a9f
		x"08", -- aa0
		x"30", -- aa1
		x"00", -- aa2
		x"0c", -- aa3
		x"12", -- aa4
		x"0e", -- aa5
		x"02", -- aa6
		x"0c", -- aa7
		x"00", -- aa8
		x"00", -- aa9
		x"00", -- aaa
		x"00", -- aab
		x"00", -- aac
		x"30", -- aad
		x"48", -- aae
		x"38", -- aaf
		x"08", -- ab0
		x"30", -- ab1
		x"00", -- ab2
		x"0c", -- ab3
		x"12", -- ab4
		x"1e", -- ab5
		x"12", -- ab6
		x"12", -- ab7
		x"00", -- ab8
		x"00", -- ab9
		x"00", -- aba
		x"00", -- abb
		x"00", -- abc
		x"30", -- abd
		x"48", -- abe
		x"38", -- abf
		x"08", -- ac0
		x"30", -- ac1
		x"00", -- ac2
		x"1c", -- ac3
		x"12", -- ac4
		x"1c", -- ac5
		x"12", -- ac6
		x"1c", -- ac7
		x"00", -- ac8
		x"00", -- ac9
		x"00", -- aca
		x"00", -- acb
		x"00", -- acc
		x"30", -- acd
		x"48", -- ace
		x"38", -- acf
		x"08", -- ad0
		x"30", -- ad1
		x"00", -- ad2
		x"0e", -- ad3
		x"10", -- ad4
		x"10", -- ad5
		x"10", -- ad6
		x"0e", -- ad7
		x"00", -- ad8
		x"00", -- ad9
		x"00", -- ada
		x"00", -- adb
		x"00", -- adc
		x"30", -- add
		x"48", -- ade
		x"38", -- adf
		x"08", -- ae0
		x"30", -- ae1
		x"00", -- ae2
		x"1c", -- ae3
		x"12", -- ae4
		x"12", -- ae5
		x"12", -- ae6
		x"1c", -- ae7
		x"00", -- ae8
		x"00", -- ae9
		x"00", -- aea
		x"00", -- aeb
		x"00", -- aec
		x"30", -- aed
		x"48", -- aee
		x"38", -- aef
		x"08", -- af0
		x"30", -- af1
		x"00", -- af2
		x"1e", -- af3
		x"10", -- af4
		x"1c", -- af5
		x"10", -- af6
		x"1e", -- af7
		x"00", -- af8
		x"00", -- af9
		x"00", -- afa
		x"00", -- afb
		x"00", -- afc
		x"30", -- afd
		x"48", -- afe
		x"38", -- aff
		x"08", -- b00
		x"30", -- b01
		x"00", -- b02
		x"1e", -- b03
		x"10", -- b04
		x"1c", -- b05
		x"10", -- b06
		x"10", -- b07
		x"00", -- b08
		x"00", -- b09
		x"00", -- b0a
		x"00", -- b0b
		x"00", -- b0c
		x"00", -- b0d
		x"00", -- b0e
		x"00", -- b0f
		x"00", -- b10
		x"00", -- b11
		x"00", -- b12
		x"00", -- b13
		x"00", -- b14
		x"00", -- b15
		x"00", -- b16
		x"00", -- b17
		x"00", -- b18
		x"00", -- b19
		x"00", -- b1a
		x"00", -- b1b
		x"10", -- b1c
		x"08", -- b1d
		x"00", -- b1e
		x"3c", -- b1f
		x"42", -- b20
		x"42", -- b21
		x"42", -- b22
		x"7e", -- b23
		x"42", -- b24
		x"42", -- b25
		x"42", -- b26
		x"42", -- b27
		x"00", -- b28
		x"00", -- b29
		x"00", -- b2a
		x"00", -- b2b
		x"10", -- b2c
		x"28", -- b2d
		x"00", -- b2e
		x"3c", -- b2f
		x"42", -- b30
		x"42", -- b31
		x"42", -- b32
		x"7e", -- b33
		x"42", -- b34
		x"42", -- b35
		x"42", -- b36
		x"42", -- b37
		x"00", -- b38
		x"00", -- b39
		x"00", -- b3a
		x"00", -- b3b
		x"10", -- b3c
		x"08", -- b3d
		x"00", -- b3e
		x"7e", -- b3f
		x"40", -- b40
		x"40", -- b41
		x"40", -- b42
		x"78", -- b43
		x"40", -- b44
		x"40", -- b45
		x"40", -- b46
		x"7e", -- b47
		x"00", -- b48
		x"00", -- b49
		x"00", -- b4a
		x"00", -- b4b
		x"10", -- b4c
		x"28", -- b4d
		x"00", -- b4e
		x"7e", -- b4f
		x"40", -- b50
		x"40", -- b51
		x"40", -- b52
		x"78", -- b53
		x"40", -- b54
		x"40", -- b55
		x"40", -- b56
		x"7e", -- b57
		x"00", -- b58
		x"00", -- b59
		x"00", -- b5a
		x"00", -- b5b
		x"00", -- b5c
		x"28", -- b5d
		x"00", -- b5e
		x"7e", -- b5f
		x"40", -- b60
		x"40", -- b61
		x"40", -- b62
		x"78", -- b63
		x"40", -- b64
		x"40", -- b65
		x"40", -- b66
		x"7e", -- b67
		x"00", -- b68
		x"00", -- b69
		x"00", -- b6a
		x"00", -- b6b
		x"10", -- b6c
		x"28", -- b6d
		x"00", -- b6e
		x"38", -- b6f
		x"10", -- b70
		x"10", -- b71
		x"10", -- b72
		x"10", -- b73
		x"10", -- b74
		x"10", -- b75
		x"10", -- b76
		x"38", -- b77
		x"00", -- b78
		x"00", -- b79
		x"00", -- b7a
		x"00", -- b7b
		x"00", -- b7c
		x"28", -- b7d
		x"00", -- b7e
		x"38", -- b7f
		x"10", -- b80
		x"10", -- b81
		x"10", -- b82
		x"10", -- b83
		x"10", -- b84
		x"10", -- b85
		x"10", -- b86
		x"38", -- b87
		x"00", -- b88
		x"00", -- b89
		x"00", -- b8a
		x"00", -- b8b
		x"08", -- b8c
		x"10", -- b8d
		x"00", -- b8e
		x"00", -- b8f
		x"00", -- b90
		x"00", -- b91
		x"00", -- b92
		x"00", -- b93
		x"00", -- b94
		x"00", -- b95
		x"00", -- b96
		x"00", -- b97
		x"00", -- b98
		x"00", -- b99
		x"00", -- b9a
		x"00", -- b9b
		x"10", -- b9c
		x"08", -- b9d
		x"00", -- b9e
		x"00", -- b9f
		x"00", -- ba0
		x"00", -- ba1
		x"00", -- ba2
		x"00", -- ba3
		x"00", -- ba4
		x"00", -- ba5
		x"00", -- ba6
		x"00", -- ba7
		x"00", -- ba8
		x"00", -- ba9
		x"00", -- baa
		x"00", -- bab
		x"10", -- bac
		x"28", -- bad
		x"00", -- bae
		x"00", -- baf
		x"00", -- bb0
		x"00", -- bb1
		x"00", -- bb2
		x"00", -- bb3
		x"00", -- bb4
		x"00", -- bb5
		x"00", -- bb6
		x"00", -- bb7
		x"00", -- bb8
		x"00", -- bb9
		x"00", -- bba
		x"00", -- bbb
		x"00", -- bbc
		x"28", -- bbd
		x"00", -- bbe
		x"00", -- bbf
		x"00", -- bc0
		x"00", -- bc1
		x"00", -- bc2
		x"00", -- bc3
		x"00", -- bc4
		x"00", -- bc5
		x"00", -- bc6
		x"00", -- bc7
		x"00", -- bc8
		x"00", -- bc9
		x"00", -- bca
		x"00", -- bcb
		x"32", -- bcc
		x"4c", -- bcd
		x"00", -- bce
		x"00", -- bcf
		x"00", -- bd0
		x"00", -- bd1
		x"00", -- bd2
		x"00", -- bd3
		x"00", -- bd4
		x"00", -- bd5
		x"00", -- bd6
		x"00", -- bd7
		x"00", -- bd8
		x"00", -- bd9
		x"00", -- bda
		x"00", -- bdb
		x"10", -- bdc
		x"08", -- bdd
		x"00", -- bde
		x"42", -- bdf
		x"42", -- be0
		x"42", -- be1
		x"42", -- be2
		x"42", -- be3
		x"42", -- be4
		x"42", -- be5
		x"42", -- be6
		x"3c", -- be7
		x"00", -- be8
		x"00", -- be9
		x"00", -- bea
		x"00", -- beb
		x"10", -- bec
		x"28", -- bed
		x"00", -- bee
		x"42", -- bef
		x"42", -- bf0
		x"42", -- bf1
		x"42", -- bf2
		x"42", -- bf3
		x"42", -- bf4
		x"42", -- bf5
		x"42", -- bf6
		x"3c", -- bf7
		x"00", -- bf8
		x"00", -- bf9
		x"00", -- bfa
		x"00", -- bfb
		x"00", -- bfc
		x"00", -- bfd
		x"0c", -- bfe
		x"12", -- bff
		x"10", -- c00
		x"3c", -- c01
		x"10", -- c02
		x"3c", -- c03
		x"10", -- c04
		x"10", -- c05
		x"51", -- c06
		x"3e", -- c07
		x"00", -- c08
		x"00", -- c09
		x"00", -- c0a
		x"00", -- c0b
		x"00", -- c0c
		x"ff", -- c0d
		x"00", -- c0e
		x"00", -- c0f
		x"00", -- c10
		x"00", -- c11
		x"00", -- c12
		x"00", -- c13
		x"00", -- c14
		x"00", -- c15
		x"00", -- c16
		x"00", -- c17
		x"00", -- c18
		x"00", -- c19
		x"00", -- c1a
		x"00", -- c1b
		x"08", -- c1c
		x"10", -- c1d
		x"00", -- c1e
		x"82", -- c1f
		x"82", -- c20
		x"44", -- c21
		x"28", -- c22
		x"10", -- c23
		x"10", -- c24
		x"10", -- c25
		x"10", -- c26
		x"10", -- c27
		x"00", -- c28
		x"00", -- c29
		x"00", -- c2a
		x"00", -- c2b
		x"08", -- c2c
		x"10", -- c2d
		x"00", -- c2e
		x"00", -- c2f
		x"00", -- c30
		x"00", -- c31
		x"42", -- c32
		x"42", -- c33
		x"42", -- c34
		x"42", -- c35
		x"42", -- c36
		x"3e", -- c37
		x"02", -- c38
		x"02", -- c39
		x"3c", -- c3a
		x"00", -- c3b
		x"00", -- c3c
		x"00", -- c3d
		x"18", -- c3e
		x"24", -- c3f
		x"24", -- c40
		x"18", -- c41
		x"00", -- c42
		x"00", -- c43
		x"00", -- c44
		x"00", -- c45
		x"00", -- c46
		x"00", -- c47
		x"00", -- c48
		x"00", -- c49
		x"00", -- c4a
		x"00", -- c4b
		x"00", -- c4c
		x"00", -- c4d
		x"3c", -- c4e
		x"42", -- c4f
		x"40", -- c50
		x"40", -- c51
		x"40", -- c52
		x"40", -- c53
		x"40", -- c54
		x"40", -- c55
		x"42", -- c56
		x"3c", -- c57
		x"10", -- c58
		x"08", -- c59
		x"10", -- c5a
		x"00", -- c5b
		x"00", -- c5c
		x"00", -- c5d
		x"00", -- c5e
		x"00", -- c5f
		x"00", -- c60
		x"00", -- c61
		x"3c", -- c62
		x"42", -- c63
		x"40", -- c64
		x"40", -- c65
		x"42", -- c66
		x"3c", -- c67
		x"10", -- c68
		x"08", -- c69
		x"10", -- c6a
		x"00", -- c6b
		x"32", -- c6c
		x"4c", -- c6d
		x"00", -- c6e
		x"42", -- c6f
		x"62", -- c70
		x"52", -- c71
		x"52", -- c72
		x"4a", -- c73
		x"4a", -- c74
		x"46", -- c75
		x"42", -- c76
		x"42", -- c77
		x"00", -- c78
		x"00", -- c79
		x"00", -- c7a
		x"00", -- c7b
		x"32", -- c7c
		x"4c", -- c7d
		x"00", -- c7e
		x"00", -- c7f
		x"00", -- c80
		x"00", -- c81
		x"5c", -- c82
		x"62", -- c83
		x"42", -- c84
		x"42", -- c85
		x"42", -- c86
		x"42", -- c87
		x"00", -- c88
		x"00", -- c89
		x"00", -- c8a
		x"00", -- c8b
		x"00", -- c8c
		x"00", -- c8d
		x"10", -- c8e
		x"00", -- c8f
		x"10", -- c90
		x"10", -- c91
		x"10", -- c92
		x"10", -- c93
		x"10", -- c94
		x"10", -- c95
		x"10", -- c96
		x"10", -- c97
		x"00", -- c98
		x"00", -- c99
		x"00", -- c9a
		x"00", -- c9b
		x"00", -- c9c
		x"00", -- c9d
		x"10", -- c9e
		x"00", -- c9f
		x"10", -- ca0
		x"10", -- ca1
		x"10", -- ca2
		x"20", -- ca3
		x"40", -- ca4
		x"40", -- ca5
		x"42", -- ca6
		x"3c", -- ca7
		x"00", -- ca8
		x"00", -- ca9
		x"00", -- caa
		x"00", -- cab
		x"00", -- cac
		x"00", -- cad
		x"00", -- cae
		x"00", -- caf
		x"00", -- cb0
		x"42", -- cb1
		x"3c", -- cb2
		x"24", -- cb3
		x"24", -- cb4
		x"24", -- cb5
		x"3c", -- cb6
		x"42", -- cb7
		x"00", -- cb8
		x"00", -- cb9
		x"00", -- cba
		x"00", -- cbb
		x"00", -- cbc
		x"00", -- cbd
		x"0c", -- cbe
		x"12", -- cbf
		x"10", -- cc0
		x"10", -- cc1
		x"3c", -- cc2
		x"10", -- cc3
		x"10", -- cc4
		x"10", -- cc5
		x"51", -- cc6
		x"3e", -- cc7
		x"00", -- cc8
		x"00", -- cc9
		x"00", -- cca
		x"00", -- ccb
		x"00", -- ccc
		x"00", -- ccd
		x"82", -- cce
		x"44", -- ccf
		x"28", -- cd0
		x"10", -- cd1
		x"7c", -- cd2
		x"10", -- cd3
		x"7c", -- cd4
		x"10", -- cd5
		x"10", -- cd6
		x"10", -- cd7
		x"00", -- cd8
		x"00", -- cd9
		x"00", -- cda
		x"00", -- cdb
		x"00", -- cdc
		x"00", -- cdd
		x"18", -- cde
		x"24", -- cdf
		x"10", -- ce0
		x"18", -- ce1
		x"24", -- ce2
		x"24", -- ce3
		x"18", -- ce4
		x"08", -- ce5
		x"24", -- ce6
		x"18", -- ce7
		x"00", -- ce8
		x"00", -- ce9
		x"00", -- cea
		x"00", -- ceb
		x"00", -- cec
		x"00", -- ced
		x"06", -- cee
		x"08", -- cef
		x"10", -- cf0
		x"10", -- cf1
		x"7c", -- cf2
		x"10", -- cf3
		x"10", -- cf4
		x"10", -- cf5
		x"20", -- cf6
		x"c0", -- cf7
		x"00", -- cf8
		x"00", -- cf9
		x"00", -- cfa
		x"00", -- cfb
		x"00", -- cfc
		x"00", -- cfd
		x"00", -- cfe
		x"00", -- cff
		x"10", -- d00
		x"38", -- d01
		x"54", -- d02
		x"50", -- d03
		x"50", -- d04
		x"54", -- d05
		x"38", -- d06
		x"10", -- d07
		x"00", -- d08
		x"00", -- d09
		x"00", -- d0a
		x"00", -- d0b
		x"10", -- d0c
		x"28", -- d0d
		x"00", -- d0e
		x"00", -- d0f
		x"00", -- d10
		x"00", -- d11
		x"3c", -- d12
		x"02", -- d13
		x"3e", -- d14
		x"42", -- d15
		x"42", -- d16
		x"3e", -- d17
		x"00", -- d18
		x"00", -- d19
		x"00", -- d1a
		x"00", -- d1b
		x"10", -- d1c
		x"28", -- d1d
		x"00", -- d1e
		x"00", -- d1f
		x"00", -- d20
		x"00", -- d21
		x"3c", -- d22
		x"42", -- d23
		x"7e", -- d24
		x"40", -- d25
		x"40", -- d26
		x"3e", -- d27
		x"00", -- d28
		x"00", -- d29
		x"00", -- d2a
		x"00", -- d2b
		x"10", -- d2c
		x"28", -- d2d
		x"00", -- d2e
		x"00", -- d2f
		x"00", -- d30
		x"00", -- d31
		x"3c", -- d32
		x"42", -- d33
		x"42", -- d34
		x"42", -- d35
		x"42", -- d36
		x"3c", -- d37
		x"00", -- d38
		x"00", -- d39
		x"00", -- d3a
		x"00", -- d3b
		x"10", -- d3c
		x"28", -- d3d
		x"00", -- d3e
		x"00", -- d3f
		x"00", -- d40
		x"00", -- d41
		x"42", -- d42
		x"42", -- d43
		x"42", -- d44
		x"42", -- d45
		x"42", -- d46
		x"3e", -- d47
		x"00", -- d48
		x"00", -- d49
		x"00", -- d4a
		x"00", -- d4b
		x"08", -- d4c
		x"10", -- d4d
		x"00", -- d4e
		x"00", -- d4f
		x"00", -- d50
		x"00", -- d51
		x"3c", -- d52
		x"02", -- d53
		x"3e", -- d54
		x"42", -- d55
		x"42", -- d56
		x"3e", -- d57
		x"00", -- d58
		x"00", -- d59
		x"00", -- d5a
		x"00", -- d5b
		x"08", -- d5c
		x"10", -- d5d
		x"00", -- d5e
		x"00", -- d5f
		x"00", -- d60
		x"00", -- d61
		x"3c", -- d62
		x"42", -- d63
		x"7e", -- d64
		x"40", -- d65
		x"40", -- d66
		x"3e", -- d67
		x"00", -- d68
		x"00", -- d69
		x"00", -- d6a
		x"00", -- d6b
		x"08", -- d6c
		x"10", -- d6d
		x"00", -- d6e
		x"00", -- d6f
		x"00", -- d70
		x"00", -- d71
		x"3c", -- d72
		x"42", -- d73
		x"42", -- d74
		x"42", -- d75
		x"42", -- d76
		x"3c", -- d77
		x"00", -- d78
		x"00", -- d79
		x"00", -- d7a
		x"00", -- d7b
		x"08", -- d7c
		x"10", -- d7d
		x"00", -- d7e
		x"00", -- d7f
		x"00", -- d80
		x"00", -- d81
		x"42", -- d82
		x"42", -- d83
		x"42", -- d84
		x"42", -- d85
		x"42", -- d86
		x"3e", -- d87
		x"00", -- d88
		x"00", -- d89
		x"00", -- d8a
		x"00", -- d8b
		x"10", -- d8c
		x"08", -- d8d
		x"00", -- d8e
		x"00", -- d8f
		x"00", -- d90
		x"00", -- d91
		x"3c", -- d92
		x"02", -- d93
		x"3e", -- d94
		x"42", -- d95
		x"42", -- d96
		x"3e", -- d97
		x"00", -- d98
		x"00", -- d99
		x"00", -- d9a
		x"00", -- d9b
		x"10", -- d9c
		x"08", -- d9d
		x"00", -- d9e
		x"00", -- d9f
		x"00", -- da0
		x"00", -- da1
		x"3c", -- da2
		x"42", -- da3
		x"7e", -- da4
		x"40", -- da5
		x"40", -- da6
		x"3e", -- da7
		x"00", -- da8
		x"00", -- da9
		x"00", -- daa
		x"00", -- dab
		x"10", -- dac
		x"08", -- dad
		x"00", -- dae
		x"00", -- daf
		x"00", -- db0
		x"00", -- db1
		x"3c", -- db2
		x"42", -- db3
		x"42", -- db4
		x"42", -- db5
		x"42", -- db6
		x"3c", -- db7
		x"00", -- db8
		x"00", -- db9
		x"00", -- dba
		x"00", -- dbb
		x"10", -- dbc
		x"08", -- dbd
		x"00", -- dbe
		x"00", -- dbf
		x"00", -- dc0
		x"00", -- dc1
		x"42", -- dc2
		x"42", -- dc3
		x"42", -- dc4
		x"42", -- dc5
		x"42", -- dc6
		x"3e", -- dc7
		x"00", -- dc8
		x"00", -- dc9
		x"00", -- dca
		x"00", -- dcb
		x"00", -- dcc
		x"28", -- dcd
		x"00", -- dce
		x"00", -- dcf
		x"00", -- dd0
		x"00", -- dd1
		x"3c", -- dd2
		x"02", -- dd3
		x"3e", -- dd4
		x"42", -- dd5
		x"42", -- dd6
		x"3e", -- dd7
		x"00", -- dd8
		x"00", -- dd9
		x"00", -- dda
		x"00", -- ddb
		x"00", -- ddc
		x"28", -- ddd
		x"00", -- dde
		x"00", -- ddf
		x"00", -- de0
		x"00", -- de1
		x"3c", -- de2
		x"42", -- de3
		x"7e", -- de4
		x"40", -- de5
		x"40", -- de6
		x"3e", -- de7
		x"00", -- de8
		x"00", -- de9
		x"00", -- dea
		x"00", -- deb
		x"00", -- dec
		x"28", -- ded
		x"00", -- dee
		x"00", -- def
		x"00", -- df0
		x"00", -- df1
		x"3c", -- df2
		x"42", -- df3
		x"42", -- df4
		x"42", -- df5
		x"42", -- df6
		x"3c", -- df7
		x"00", -- df8
		x"00", -- df9
		x"00", -- dfa
		x"00", -- dfb
		x"00", -- dfc
		x"28", -- dfd
		x"00", -- dfe
		x"00", -- dff
		x"00", -- e00
		x"00", -- e01
		x"42", -- e02
		x"42", -- e03
		x"42", -- e04
		x"42", -- e05
		x"42", -- e06
		x"3e", -- e07
		x"00", -- e08
		x"00", -- e09
		x"00", -- e0a
		x"00", -- e0b
		x"18", -- e0c
		x"18", -- e0d
		x"00", -- e0e
		x"3c", -- e0f
		x"42", -- e10
		x"42", -- e11
		x"42", -- e12
		x"7e", -- e13
		x"42", -- e14
		x"42", -- e15
		x"42", -- e16
		x"42", -- e17
		x"00", -- e18
		x"00", -- e19
		x"00", -- e1a
		x"00", -- e1b
		x"10", -- e1c
		x"28", -- e1d
		x"00", -- e1e
		x"00", -- e1f
		x"00", -- e20
		x"00", -- e21
		x"30", -- e22
		x"10", -- e23
		x"10", -- e24
		x"10", -- e25
		x"10", -- e26
		x"38", -- e27
		x"00", -- e28
		x"00", -- e29
		x"00", -- e2a
		x"00", -- e2b
		x"00", -- e2c
		x"00", -- e2d
		x"3d", -- e2e
		x"42", -- e2f
		x"46", -- e30
		x"4a", -- e31
		x"4a", -- e32
		x"52", -- e33
		x"52", -- e34
		x"62", -- e35
		x"42", -- e36
		x"bc", -- e37
		x"00", -- e38
		x"00", -- e39
		x"00", -- e3a
		x"00", -- e3b
		x"00", -- e3c
		x"00", -- e3d
		x"3f", -- e3e
		x"48", -- e3f
		x"48", -- e40
		x"48", -- e41
		x"7e", -- e42
		x"48", -- e43
		x"48", -- e44
		x"48", -- e45
		x"48", -- e46
		x"4f", -- e47
		x"00", -- e48
		x"00", -- e49
		x"00", -- e4a
		x"00", -- e4b
		x"18", -- e4c
		x"18", -- e4d
		x"00", -- e4e
		x"00", -- e4f
		x"00", -- e50
		x"00", -- e51
		x"3c", -- e52
		x"02", -- e53
		x"3e", -- e54
		x"42", -- e55
		x"42", -- e56
		x"3e", -- e57
		x"00", -- e58
		x"00", -- e59
		x"00", -- e5a
		x"00", -- e5b
		x"08", -- e5c
		x"10", -- e5d
		x"00", -- e5e
		x"00", -- e5f
		x"00", -- e60
		x"00", -- e61
		x"30", -- e62
		x"10", -- e63
		x"10", -- e64
		x"10", -- e65
		x"10", -- e66
		x"38", -- e67
		x"00", -- e68
		x"00", -- e69
		x"00", -- e6a
		x"00", -- e6b
		x"00", -- e6c
		x"00", -- e6d
		x"00", -- e6e
		x"00", -- e6f
		x"00", -- e70
		x"00", -- e71
		x"3d", -- e72
		x"42", -- e73
		x"4e", -- e74
		x"72", -- e75
		x"42", -- e76
		x"bc", -- e77
		x"00", -- e78
		x"00", -- e79
		x"00", -- e7a
		x"00", -- e7b
		x"00", -- e7c
		x"00", -- e7d
		x"00", -- e7e
		x"00", -- e7f
		x"00", -- e80
		x"00", -- e81
		x"36", -- e82
		x"09", -- e83
		x"3f", -- e84
		x"48", -- e85
		x"49", -- e86
		x"36", -- e87
		x"00", -- e88
		x"00", -- e89
		x"00", -- e8a
		x"00", -- e8b
		x"00", -- e8c
		x"28", -- e8d
		x"00", -- e8e
		x"3c", -- e8f
		x"42", -- e90
		x"42", -- e91
		x"42", -- e92
		x"7e", -- e93
		x"42", -- e94
		x"42", -- e95
		x"42", -- e96
		x"42", -- e97
		x"00", -- e98
		x"00", -- e99
		x"00", -- e9a
		x"00", -- e9b
		x"10", -- e9c
		x"08", -- e9d
		x"00", -- e9e
		x"00", -- e9f
		x"00", -- ea0
		x"00", -- ea1
		x"30", -- ea2
		x"10", -- ea3
		x"10", -- ea4
		x"10", -- ea5
		x"10", -- ea6
		x"38", -- ea7
		x"00", -- ea8
		x"00", -- ea9
		x"00", -- eaa
		x"00", -- eab
		x"00", -- eac
		x"28", -- ead
		x"00", -- eae
		x"3c", -- eaf
		x"42", -- eb0
		x"42", -- eb1
		x"42", -- eb2
		x"42", -- eb3
		x"42", -- eb4
		x"42", -- eb5
		x"42", -- eb6
		x"3c", -- eb7
		x"00", -- eb8
		x"00", -- eb9
		x"00", -- eba
		x"00", -- ebb
		x"00", -- ebc
		x"28", -- ebd
		x"00", -- ebe
		x"42", -- ebf
		x"42", -- ec0
		x"42", -- ec1
		x"42", -- ec2
		x"42", -- ec3
		x"42", -- ec4
		x"42", -- ec5
		x"42", -- ec6
		x"3c", -- ec7
		x"00", -- ec8
		x"00", -- ec9
		x"00", -- eca
		x"00", -- ecb
		x"08", -- ecc
		x"10", -- ecd
		x"00", -- ece
		x"7e", -- ecf
		x"40", -- ed0
		x"40", -- ed1
		x"40", -- ed2
		x"78", -- ed3
		x"40", -- ed4
		x"40", -- ed5
		x"40", -- ed6
		x"7e", -- ed7
		x"00", -- ed8
		x"00", -- ed9
		x"00", -- eda
		x"00", -- edb
		x"00", -- edc
		x"28", -- edd
		x"00", -- ede
		x"00", -- edf
		x"00", -- ee0
		x"00", -- ee1
		x"30", -- ee2
		x"10", -- ee3
		x"10", -- ee4
		x"10", -- ee5
		x"10", -- ee6
		x"38", -- ee7
		x"00", -- ee8
		x"00", -- ee9
		x"00", -- eea
		x"00", -- eeb
		x"00", -- eec
		x"00", -- eed
		x"18", -- eee
		x"24", -- eef
		x"44", -- ef0
		x"48", -- ef1
		x"70", -- ef2
		x"48", -- ef3
		x"44", -- ef4
		x"44", -- ef5
		x"64", -- ef6
		x"58", -- ef7
		x"00", -- ef8
		x"00", -- ef9
		x"00", -- efa
		x"00", -- efb
		x"10", -- efc
		x"28", -- efd
		x"00", -- efe
		x"3c", -- eff
		x"42", -- f00
		x"42", -- f01
		x"42", -- f02
		x"42", -- f03
		x"42", -- f04
		x"42", -- f05
		x"42", -- f06
		x"3c", -- f07
		x"00", -- f08
		x"00", -- f09
		x"00", -- f0a
		x"00", -- f0b
		x"08", -- f0c
		x"10", -- f0d
		x"00", -- f0e
		x"3c", -- f0f
		x"42", -- f10
		x"42", -- f11
		x"42", -- f12
		x"7e", -- f13
		x"42", -- f14
		x"42", -- f15
		x"42", -- f16
		x"42", -- f17
		x"00", -- f18
		x"00", -- f19
		x"00", -- f1a
		x"00", -- f1b
		x"32", -- f1c
		x"4c", -- f1d
		x"00", -- f1e
		x"3c", -- f1f
		x"42", -- f20
		x"42", -- f21
		x"42", -- f22
		x"7e", -- f23
		x"42", -- f24
		x"42", -- f25
		x"42", -- f26
		x"42", -- f27
		x"00", -- f28
		x"00", -- f29
		x"00", -- f2a
		x"00", -- f2b
		x"32", -- f2c
		x"4c", -- f2d
		x"00", -- f2e
		x"00", -- f2f
		x"00", -- f30
		x"00", -- f31
		x"3c", -- f32
		x"02", -- f33
		x"3e", -- f34
		x"42", -- f35
		x"42", -- f36
		x"3e", -- f37
		x"00", -- f38
		x"00", -- f39
		x"00", -- f3a
		x"00", -- f3b
		x"00", -- f3c
		x"00", -- f3d
		x"7c", -- f3e
		x"42", -- f3f
		x"42", -- f40
		x"42", -- f41
		x"e2", -- f42
		x"42", -- f43
		x"42", -- f44
		x"42", -- f45
		x"42", -- f46
		x"7c", -- f47
		x"00", -- f48
		x"00", -- f49
		x"00", -- f4a
		x"00", -- f4b
		x"00", -- f4c
		x"00", -- f4d
		x"00", -- f4e
		x"04", -- f4f
		x"0e", -- f50
		x"04", -- f51
		x"3c", -- f52
		x"44", -- f53
		x"44", -- f54
		x"44", -- f55
		x"44", -- f56
		x"38", -- f57
		x"00", -- f58
		x"00", -- f59
		x"00", -- f5a
		x"00", -- f5b
		x"08", -- f5c
		x"10", -- f5d
		x"00", -- f5e
		x"38", -- f5f
		x"10", -- f60
		x"10", -- f61
		x"10", -- f62
		x"10", -- f63
		x"10", -- f64
		x"10", -- f65
		x"10", -- f66
		x"38", -- f67
		x"00", -- f68
		x"00", -- f69
		x"00", -- f6a
		x"00", -- f6b
		x"10", -- f6c
		x"08", -- f6d
		x"00", -- f6e
		x"38", -- f6f
		x"10", -- f70
		x"10", -- f71
		x"10", -- f72
		x"10", -- f73
		x"10", -- f74
		x"10", -- f75
		x"10", -- f76
		x"38", -- f77
		x"00", -- f78
		x"00", -- f79
		x"00", -- f7a
		x"00", -- f7b
		x"08", -- f7c
		x"10", -- f7d
		x"00", -- f7e
		x"3c", -- f7f
		x"42", -- f80
		x"42", -- f81
		x"42", -- f82
		x"42", -- f83
		x"42", -- f84
		x"42", -- f85
		x"42", -- f86
		x"3c", -- f87
		x"00", -- f88
		x"00", -- f89
		x"00", -- f8a
		x"00", -- f8b
		x"10", -- f8c
		x"08", -- f8d
		x"00", -- f8e
		x"3c", -- f8f
		x"42", -- f90
		x"42", -- f91
		x"42", -- f92
		x"42", -- f93
		x"42", -- f94
		x"42", -- f95
		x"42", -- f96
		x"3c", -- f97
		x"00", -- f98
		x"00", -- f99
		x"00", -- f9a
		x"00", -- f9b
		x"32", -- f9c
		x"4c", -- f9d
		x"00", -- f9e
		x"3c", -- f9f
		x"42", -- fa0
		x"42", -- fa1
		x"42", -- fa2
		x"42", -- fa3
		x"42", -- fa4
		x"42", -- fa5
		x"42", -- fa6
		x"3c", -- fa7
		x"00", -- fa8
		x"00", -- fa9
		x"00", -- faa
		x"00", -- fab
		x"32", -- fac
		x"4c", -- fad
		x"00", -- fae
		x"00", -- faf
		x"00", -- fb0
		x"00", -- fb1
		x"3c", -- fb2
		x"42", -- fb3
		x"42", -- fb4
		x"42", -- fb5
		x"42", -- fb6
		x"3c", -- fb7
		x"00", -- fb8
		x"00", -- fb9
		x"00", -- fba
		x"00", -- fbb
		x"28", -- fbc
		x"10", -- fbd
		x"00", -- fbe
		x"3c", -- fbf
		x"42", -- fc0
		x"40", -- fc1
		x"40", -- fc2
		x"3c", -- fc3
		x"02", -- fc4
		x"02", -- fc5
		x"42", -- fc6
		x"3c", -- fc7
		x"00", -- fc8
		x"00", -- fc9
		x"00", -- fca
		x"00", -- fcb
		x"28", -- fcc
		x"10", -- fcd
		x"00", -- fce
		x"00", -- fcf
		x"00", -- fd0
		x"00", -- fd1
		x"3c", -- fd2
		x"40", -- fd3
		x"3c", -- fd4
		x"02", -- fd5
		x"42", -- fd6
		x"3c", -- fd7
		x"00", -- fd8
		x"00", -- fd9
		x"00", -- fda
		x"00", -- fdb
		x"08", -- fdc
		x"10", -- fdd
		x"00", -- fde
		x"42", -- fdf
		x"42", -- fe0
		x"42", -- fe1
		x"42", -- fe2
		x"42", -- fe3
		x"42", -- fe4
		x"42", -- fe5
		x"42", -- fe6
		x"3c", -- fe7
		x"00", -- fe8
		x"00", -- fe9
		x"00", -- fea
		x"00", -- feb
		x"00", -- fec
		x"28", -- fed
		x"00", -- fee
		x"82", -- fef
		x"82", -- ff0
		x"44", -- ff1
		x"28", -- ff2
		x"10", -- ff3
		x"10", -- ff4
		x"10", -- ff5
		x"10", -- ff6
		x"10", -- ff7
		x"00", -- ff8
		x"00", -- ff9
		x"00", -- ffa
		x"00", -- ffb
		x"00", -- ffc
		x"28", -- ffd
		x"00", -- ffe
		x"00", -- fff
		x"00", -- 1000
		x"00", -- 1001
		x"42", -- 1002
		x"42", -- 1003
		x"42", -- 1004
		x"42", -- 1005
		x"42", -- 1006
		x"3e", -- 1007
		x"02", -- 1008
		x"02", -- 1009
		x"3c", -- 100a
		x"00", -- 100b
		x"00", -- 100c
		x"00", -- 100d
		x"38", -- 100e
		x"10", -- 100f
		x"10", -- 1010
		x"1c", -- 1011
		x"12", -- 1012
		x"12", -- 1013
		x"1c", -- 1014
		x"10", -- 1015
		x"10", -- 1016
		x"38", -- 1017
		x"00", -- 1018
		x"00", -- 1019
		x"00", -- 101a
		x"00", -- 101b
		x"00", -- 101c
		x"00", -- 101d
		x"00", -- 101e
		x"00", -- 101f
		x"10", -- 1020
		x"10", -- 1021
		x"1c", -- 1022
		x"12", -- 1023
		x"12", -- 1024
		x"1c", -- 1025
		x"10", -- 1026
		x"10", -- 1027
		x"00", -- 1028
		x"00", -- 1029
		x"00", -- 102a
		x"00", -- 102b
		x"00", -- 102c
		x"00", -- 102d
		x"00", -- 102e
		x"00", -- 102f
		x"00", -- 1030
		x"00", -- 1031
		x"30", -- 1032
		x"30", -- 1033
		x"00", -- 1034
		x"00", -- 1035
		x"00", -- 1036
		x"00", -- 1037
		x"00", -- 1038
		x"00", -- 1039
		x"00", -- 103a
		x"00", -- 103b
		x"00", -- 103c
		x"00", -- 103d
		x"00", -- 103e
		x"00", -- 103f
		x"00", -- 1040
		x"00", -- 1041
		x"44", -- 1042
		x"44", -- 1043
		x"44", -- 1044
		x"44", -- 1045
		x"64", -- 1046
		x"5a", -- 1047
		x"40", -- 1048
		x"40", -- 1049
		x"00", -- 104a
		x"00", -- 104b
		x"00", -- 104c
		x"00", -- 104d
		x"7e", -- 104e
		x"f4", -- 104f
		x"f4", -- 1050
		x"f4", -- 1051
		x"f4", -- 1052
		x"74", -- 1053
		x"14", -- 1054
		x"14", -- 1055
		x"14", -- 1056
		x"14", -- 1057
		x"00", -- 1058
		x"00", -- 1059
		x"00", -- 105a
		x"00", -- 105b
		x"00", -- 105c
		x"70", -- 105d
		x"20", -- 105e
		x"20", -- 105f
		x"20", -- 1060
		x"70", -- 1061
		x"00", -- 1062
		x"0c", -- 1063
		x"12", -- 1064
		x"12", -- 1065
		x"12", -- 1066
		x"0c", -- 1067
		x"00", -- 1068
		x"00", -- 1069
		x"00", -- 106a
		x"00", -- 106b
		x"00", -- 106c
		x"00", -- 106d
		x"00", -- 106e
		x"00", -- 106f
		x"00", -- 1070
		x"00", -- 1071
		x"ff", -- 1072
		x"00", -- 1073
		x"00", -- 1074
		x"00", -- 1075
		x"00", -- 1076
		x"00", -- 1077
		x"00", -- 1078
		x"00", -- 1079
		x"00", -- 107a
		x"00", -- 107b
		x"00", -- 107c
		x"20", -- 107d
		x"60", -- 107e
		x"22", -- 107f
		x"24", -- 1080
		x"28", -- 1081
		x"14", -- 1082
		x"2c", -- 1083
		x"54", -- 1084
		x"1e", -- 1085
		x"04", -- 1086
		x"0e", -- 1087
		x"00", -- 1088
		x"00", -- 1089
		x"00", -- 108a
		x"00", -- 108b
		x"00", -- 108c
		x"20", -- 108d
		x"60", -- 108e
		x"22", -- 108f
		x"24", -- 1090
		x"28", -- 1091
		x"10", -- 1092
		x"2c", -- 1093
		x"52", -- 1094
		x"04", -- 1095
		x"08", -- 1096
		x"1e", -- 1097
		x"00", -- 1098
		x"00", -- 1099
		x"00", -- 109a
		x"00", -- 109b
		x"00", -- 109c
		x"00", -- 109d
		x"3c", -- 109e
		x"02", -- 109f
		x"3e", -- 10a0
		x"42", -- 10a1
		x"3e", -- 10a2
		x"00", -- 10a3
		x"7e", -- 10a4
		x"00", -- 10a5
		x"00", -- 10a6
		x"00", -- 10a7
		x"00", -- 10a8
		x"00", -- 10a9
		x"00", -- 10aa
		x"00", -- 10ab
		x"00", -- 10ac
		x"00", -- 10ad
		x"3c", -- 10ae
		x"42", -- 10af
		x"42", -- 10b0
		x"42", -- 10b1
		x"3c", -- 10b2
		x"00", -- 10b3
		x"7e", -- 10b4
		x"00", -- 10b5
		x"00", -- 10b6
		x"00", -- 10b7
		x"00", -- 10b8
		x"00", -- 10b9
		x"00", -- 10ba
		x"00", -- 10bb
		x"00", -- 10bc
		x"00", -- 10bd
		x"09", -- 10be
		x"12", -- 10bf
		x"24", -- 10c0
		x"48", -- 10c1
		x"24", -- 10c2
		x"12", -- 10c3
		x"09", -- 10c4
		x"00", -- 10c5
		x"00", -- 10c6
		x"00", -- 10c7
		x"00", -- 10c8
		x"00", -- 10c9
		x"00", -- 10ca
		x"00", -- 10cb
		x"00", -- 10cc
		x"00", -- 10cd
		x"7e", -- 10ce
		x"7e", -- 10cf
		x"7e", -- 10d0
		x"7e", -- 10d1
		x"7e", -- 10d2
		x"7e", -- 10d3
		x"7e", -- 10d4
		x"7e", -- 10d5
		x"7e", -- 10d6
		x"00", -- 10d7
		x"00", -- 10d8
		x"00", -- 10d9
		x"00", -- 10da
		x"00", -- 10db
		x"00", -- 10dc
		x"00", -- 10dd
		x"48", -- 10de
		x"24", -- 10df
		x"12", -- 10e0
		x"09", -- 10e1
		x"12", -- 10e2
		x"24", -- 10e3
		x"48", -- 10e4
		x"00", -- 10e5
		x"00", -- 10e6
		x"00", -- 10e7
		x"00", -- 10e8
		x"00", -- 10e9
		x"00", -- 10ea
		x"00", -- 10eb
		x"00", -- 10ec
		x"00", -- 10ed
		x"00", -- 10ee
		x"10", -- 10ef
		x"10", -- 10f0
		x"7c", -- 10f1
		x"10", -- 10f2
		x"10", -- 10f3
		x"00", -- 10f4
		x"fe", -- 10f5
		x"00", -- 10f6
		x"00", -- 10f7
		x"00", -- 10f8
		x"00", -- 10f9
		x"00", -- 10fa
		x"00", -- 10fb
		x"00", -- 10fc
		x"00", -- 10fd
		x"3c", -- 10fe
		x"7e", -- 10ff
		x"5a", -- 1100
		x"56", -- 1101
		x"4e", -- 1102
		x"4e", -- 1103
		x"56", -- 1104
		x"5a", -- 1105
		x"7e", -- 1106
		x"3c", -- 1107
		x"00", -- 1108
		x"00", -- 1109
		x"00", -- 110a
		x"00", -- 110b
		x"10", -- 110c
		x"08", -- 110d
		x"01", -- 110e
		x"80", -- 110f
		x"ff", -- 1110
		x"00", -- 1111
		x"38", -- 1112
		x"40", -- 1113
		x"40", -- 1114
		x"40", -- 1115
		x"38", -- 1116
		x"00", -- 1117
		x"10", -- 1118
		x"10", -- 1119
		x"10", -- 111a
		x"10", -- 111b
		x"1e", -- 111c
		x"00", -- 111d
		x"00", -- 111e
		x"00", -- 111f
		x"00", -- 1120
		x"00", -- 1121
		x"70", -- 1122
		x"20", -- 1123
		x"20", -- 1124
		x"20", -- 1125
		x"70", -- 1126
		x"00", -- 1127
		x"22", -- 1128
		x"22", -- 1129
		x"14", -- 112a
		x"14", -- 112b
		x"08", -- 112c
		x"00", -- 112d
		x"00", -- 112e
		x"00", -- 112f
		x"00", -- 1130
		x"00", -- 1131
		x"70", -- 1132
		x"48", -- 1133
		x"70", -- 1134
		x"48", -- 1135
		x"70", -- 1136
		x"00", -- 1137
		x"0c", -- 1138
		x"10", -- 1139
		x"16", -- 113a
		x"12", -- 113b
		x"0c", -- 113c
		x"00", -- 113d
		x"00", -- 113e
		x"00", -- 113f
		x"00", -- 1140
		x"00", -- 1141
		x"70", -- 1142
		x"20", -- 1143
		x"20", -- 1144
		x"20", -- 1145
		x"70", -- 1146
		x"00", -- 1147
		x"1c", -- 1148
		x"12", -- 1149
		x"1c", -- 114a
		x"12", -- 114b
		x"1c", -- 114c
		x"00", -- 114d
		x"00", -- 114e
		x"00", -- 114f
		x"00", -- 1150
		x"00", -- 1151
		x"48", -- 1152
		x"48", -- 1153
		x"48", -- 1154
		x"48", -- 1155
		x"30", -- 1156
		x"00", -- 1157
		x"10", -- 1158
		x"10", -- 1159
		x"10", -- 115a
		x"10", -- 115b
		x"1e", -- 115c
		x"00", -- 115d
		x"ff", -- 115e
		x"00", -- 115f
		x"00", -- 1160
		x"00", -- 1161
		x"70", -- 1162
		x"20", -- 1163
		x"20", -- 1164
		x"20", -- 1165
		x"70", -- 1166
		x"00", -- 1167
		x"22", -- 1168
		x"22", -- 1169
		x"14", -- 116a
		x"14", -- 116b
		x"08", -- 116c
		x"00", -- 116d
		x"ff", -- 116e
		x"00", -- 116f
		x"00", -- 1170
		x"00", -- 1171
		x"70", -- 1172
		x"48", -- 1173
		x"70", -- 1174
		x"48", -- 1175
		x"70", -- 1176
		x"00", -- 1177
		x"0c", -- 1178
		x"10", -- 1179
		x"16", -- 117a
		x"12", -- 117b
		x"0c", -- 117c
		x"00", -- 117d
		x"ff", -- 117e
		x"00", -- 117f
		x"00", -- 1180
		x"00", -- 1181
		x"70", -- 1182
		x"20", -- 1183
		x"20", -- 1184
		x"20", -- 1185
		x"70", -- 1186
		x"00", -- 1187
		x"1c", -- 1188
		x"12", -- 1189
		x"1c", -- 118a
		x"12", -- 118b
		x"1c", -- 118c
		x"00", -- 118d
		x"ff", -- 118e
		x"00", -- 118f
		x"00", -- 1190
		x"00", -- 1191
		x"a8", -- 1192
		x"a8", -- 1193
		x"a8", -- 1194
		x"a8", -- 1195
		x"50", -- 1196
		x"00", -- 1197
		x"12", -- 1198
		x"12", -- 1199
		x"1e", -- 119a
		x"12", -- 119b
		x"12", -- 119c
		x"00", -- 119d
		x"00", -- 119e
		x"00", -- 119f
		x"00", -- 11a0
		x"00", -- 11a1
		x"70", -- 11a2
		x"48", -- 11a3
		x"70", -- 11a4
		x"50", -- 11a5
		x"48", -- 11a6
		x"00", -- 11a7
		x"1c", -- 11a8
		x"12", -- 11a9
		x"12", -- 11aa
		x"12", -- 11ab
		x"1c", -- 11ac
		x"00", -- 11ad
		x"00", -- 11ae
		x"00", -- 11af
		x"00", -- 11b0
		x"00", -- 11b1
		x"44", -- 11b2
		x"28", -- 11b3
		x"10", -- 11b4
		x"10", -- 11b5
		x"10", -- 11b6
		x"00", -- 11b7
		x"1e", -- 11b8
		x"10", -- 11b9
		x"1c", -- 11ba
		x"10", -- 11bb
		x"1e", -- 11bc
		x"00", -- 11bd
		x"00", -- 11be
		x"00", -- 11bf
		x"00", -- 11c0
		x"00", -- 11c1
		x"30", -- 11c2
		x"40", -- 11c3
		x"58", -- 11c4
		x"48", -- 11c5
		x"30", -- 11c6
		x"00", -- 11c7
		x"1c", -- 11c8
		x"12", -- 11c9
		x"1c", -- 11ca
		x"14", -- 11cb
		x"12", -- 11cc
		x"00", -- 11cd
		x"00", -- 11ce
		x"00", -- 11cf
		x"00", -- 11d0
		x"00", -- 11d1
		x"38", -- 11d2
		x"40", -- 11d3
		x"40", -- 11d4
		x"40", -- 11d5
		x"38", -- 11d6
		x"00", -- 11d7
		x"22", -- 11d8
		x"14", -- 11d9
		x"08", -- 11da
		x"08", -- 11db
		x"08", -- 11dc
		x"00", -- 11dd
		x"00", -- 11de
		x"00", -- 11df
		x"00", -- 11e0
		x"00", -- 11e1
		x"70", -- 11e2
		x"48", -- 11e3
		x"70", -- 11e4
		x"48", -- 11e5
		x"70", -- 11e6
		x"00", -- 11e7
		x"12", -- 11e8
		x"12", -- 11e9
		x"12", -- 11ea
		x"12", -- 11eb
		x"0c", -- 11ec
		x"00", -- 11ed
		x"00", -- 11ee
		x"00", -- 11ef
		x"00", -- 11f0
		x"00", -- 11f1
		x"88", -- 11f2
		x"d8", -- 11f3
		x"a8", -- 11f4
		x"88", -- 11f5
		x"88", -- 11f6
		x"00", -- 11f7
		x"0c", -- 11f8
		x"10", -- 11f9
		x"16", -- 11fa
		x"12", -- 11fb
		x"0c", -- 11fc
		x"00", -- 11fd
		x"00", -- 11fe
		x"00", -- 11ff
		x"00", -- 1200
		x"00", -- 1201
		x"70", -- 1202
		x"48", -- 1203
		x"70", -- 1204
		x"48", -- 1205
		x"70", -- 1206
		x"00", -- 1207
		x"12", -- 1208
		x"14", -- 1209
		x"18", -- 120a
		x"14", -- 120b
		x"12", -- 120c
		x"00", -- 120d
		x"00", -- 120e
		x"00", -- 120f
		x"00", -- 1210
		x"00", -- 1211
		x"30", -- 1212
		x"48", -- 1213
		x"38", -- 1214
		x"08", -- 1215
		x"30", -- 1216
		x"00", -- 1217
		x"0c", -- 1218
		x"12", -- 1219
		x"12", -- 121a
		x"12", -- 121b
		x"0c", -- 121c
		x"00", -- 121d
		x"00", -- 121e
		x"00", -- 121f
		x"00", -- 1220
		x"00", -- 1221
		x"30", -- 1222
		x"48", -- 1223
		x"38", -- 1224
		x"08", -- 1225
		x"30", -- 1226
		x"00", -- 1227
		x"04", -- 1228
		x"0c", -- 1229
		x"04", -- 122a
		x"04", -- 122b
		x"0e", -- 122c
		x"00", -- 122d
		x"00", -- 122e
		x"00", -- 122f
		x"00", -- 1230
		x"00", -- 1231
		x"30", -- 1232
		x"48", -- 1233
		x"38", -- 1234
		x"08", -- 1235
		x"30", -- 1236
		x"00", -- 1237
		x"0c", -- 1238
		x"12", -- 1239
		x"04", -- 123a
		x"08", -- 123b
		x"1e", -- 123c
		x"00", -- 123d
		x"00", -- 123e
		x"00", -- 123f
		x"00", -- 1240
		x"00", -- 1241
		x"30", -- 1242
		x"48", -- 1243
		x"38", -- 1244
		x"08", -- 1245
		x"30", -- 1246
		x"00", -- 1247
		x"1c", -- 1248
		x"02", -- 1249
		x"1c", -- 124a
		x"02", -- 124b
		x"1c", -- 124c
		x"00", -- 124d
		x"00", -- 124e
		x"00", -- 124f
		x"00", -- 1250
		x"00", -- 1251
		x"30", -- 1252
		x"48", -- 1253
		x"38", -- 1254
		x"08", -- 1255
		x"30", -- 1256
		x"00", -- 1257
		x"14", -- 1258
		x"14", -- 1259
		x"1e", -- 125a
		x"04", -- 125b
		x"04", -- 125c
		x"00", -- 125d
		x"00", -- 125e
		x"00", -- 125f
		x"00", -- 1260
		x"00", -- 1261
		x"30", -- 1262
		x"48", -- 1263
		x"38", -- 1264
		x"08", -- 1265
		x"30", -- 1266
		x"00", -- 1267
		x"1e", -- 1268
		x"10", -- 1269
		x"1c", -- 126a
		x"02", -- 126b
		x"1c", -- 126c
		x"00", -- 126d
		x"00", -- 126e
		x"00", -- 126f
		x"00", -- 1270
		x"00", -- 1271
		x"30", -- 1272
		x"48", -- 1273
		x"38", -- 1274
		x"08", -- 1275
		x"30", -- 1276
		x"00", -- 1277
		x"0c", -- 1278
		x"10", -- 1279
		x"1c", -- 127a
		x"12", -- 127b
		x"0c", -- 127c
		x"00", -- 127d
		x"00", -- 127e
		x"00", -- 127f
		x"00", -- 1280
		x"00", -- 1281
		x"30", -- 1282
		x"48", -- 1283
		x"38", -- 1284
		x"08", -- 1285
		x"30", -- 1286
		x"00", -- 1287
		x"1e", -- 1288
		x"02", -- 1289
		x"04", -- 128a
		x"08", -- 128b
		x"10", -- 128c
		x"00", -- 128d
		x"00", -- 128e
		x"00", -- 128f
		x"00", -- 1290
		x"00", -- 1291
		x"30", -- 1292
		x"48", -- 1293
		x"38", -- 1294
		x"08", -- 1295
		x"30", -- 1296
		x"00", -- 1297
		x"0c", -- 1298
		x"12", -- 1299
		x"0c", -- 129a
		x"12", -- 129b
		x"0c", -- 129c
		x"00", -- 129d
		x"00", -- 129e
		x"00", -- 129f
		x"00", -- 12a0
		x"00", -- 12a1
		x"30", -- 12a2
		x"48", -- 12a3
		x"38", -- 12a4
		x"08", -- 12a5
		x"30", -- 12a6
		x"00", -- 12a7
		x"0c", -- 12a8
		x"12", -- 12a9
		x"0e", -- 12aa
		x"02", -- 12ab
		x"0c", -- 12ac
		x"00", -- 12ad
		x"00", -- 12ae
		x"00", -- 12af
		x"00", -- 12b0
		x"00", -- 12b1
		x"30", -- 12b2
		x"48", -- 12b3
		x"38", -- 12b4
		x"08", -- 12b5
		x"30", -- 12b6
		x"00", -- 12b7
		x"0c", -- 12b8
		x"12", -- 12b9
		x"1e", -- 12ba
		x"12", -- 12bb
		x"12", -- 12bc
		x"00", -- 12bd
		x"00", -- 12be
		x"00", -- 12bf
		x"00", -- 12c0
		x"00", -- 12c1
		x"30", -- 12c2
		x"48", -- 12c3
		x"38", -- 12c4
		x"08", -- 12c5
		x"30", -- 12c6
		x"00", -- 12c7
		x"1c", -- 12c8
		x"12", -- 12c9
		x"1c", -- 12ca
		x"12", -- 12cb
		x"1c", -- 12cc
		x"00", -- 12cd
		x"00", -- 12ce
		x"00", -- 12cf
		x"00", -- 12d0
		x"00", -- 12d1
		x"30", -- 12d2
		x"48", -- 12d3
		x"38", -- 12d4
		x"08", -- 12d5
		x"30", -- 12d6
		x"00", -- 12d7
		x"0e", -- 12d8
		x"10", -- 12d9
		x"10", -- 12da
		x"10", -- 12db
		x"0e", -- 12dc
		x"00", -- 12dd
		x"00", -- 12de
		x"00", -- 12df
		x"00", -- 12e0
		x"00", -- 12e1
		x"30", -- 12e2
		x"48", -- 12e3
		x"38", -- 12e4
		x"08", -- 12e5
		x"30", -- 12e6
		x"00", -- 12e7
		x"1c", -- 12e8
		x"12", -- 12e9
		x"12", -- 12ea
		x"12", -- 12eb
		x"1c", -- 12ec
		x"00", -- 12ed
		x"00", -- 12ee
		x"00", -- 12ef
		x"00", -- 12f0
		x"00", -- 12f1
		x"30", -- 12f2
		x"48", -- 12f3
		x"38", -- 12f4
		x"08", -- 12f5
		x"30", -- 12f6
		x"00", -- 12f7
		x"1e", -- 12f8
		x"10", -- 12f9
		x"1c", -- 12fa
		x"10", -- 12fb
		x"1e", -- 12fc
		x"00", -- 12fd
		x"00", -- 12fe
		x"00", -- 12ff
		x"00", -- 1300
		x"00", -- 1301
		x"30", -- 1302
		x"48", -- 1303
		x"38", -- 1304
		x"08", -- 1305
		x"30", -- 1306
		x"00", -- 1307
		x"1e", -- 1308
		x"10", -- 1309
		x"1c", -- 130a
		x"10", -- 130b
		x"10", -- 130c
		x"00", -- 130d
		x"00", -- 130e
		x"00", -- 130f
		x"00", -- 1310
		x"00", -- 1311
		x"00", -- 1312
		x"00", -- 1313
		x"00", -- 1314
		x"00", -- 1315
		x"00", -- 1316
		x"00", -- 1317
		x"00", -- 1318
		x"00", -- 1319
		x"00", -- 131a
		x"00", -- 131b
		x"00", -- 131c
		x"00", -- 131d
		x"00", -- 131e
		x"00", -- 131f
		x"00", -- 1320
		x"00", -- 1321
		x"00", -- 1322
		x"00", -- 1323
		x"00", -- 1324
		x"00", -- 1325
		x"00", -- 1326
		x"00", -- 1327
		x"00", -- 1328
		x"00", -- 1329
		x"00", -- 132a
		x"30", -- 132b
		x"30", -- 132c
		x"00", -- 132d
		x"00", -- 132e
		x"00", -- 132f
		x"00", -- 1330
		x"00", -- 1331
		x"00", -- 1332
		x"00", -- 1333
		x"3c", -- 1334
		x"20", -- 1335
		x"20", -- 1336
		x"20", -- 1337
		x"20", -- 1338
		x"20", -- 1339
		x"20", -- 133a
		x"20", -- 133b
		x"20", -- 133c
		x"00", -- 133d
		x"00", -- 133e
		x"00", -- 133f
		x"00", -- 1340
		x"00", -- 1341
		x"00", -- 1342
		x"00", -- 1343
		x"04", -- 1344
		x"04", -- 1345
		x"04", -- 1346
		x"04", -- 1347
		x"04", -- 1348
		x"04", -- 1349
		x"04", -- 134a
		x"04", -- 134b
		x"3c", -- 134c
		x"00", -- 134d
		x"00", -- 134e
		x"00", -- 134f
		x"00", -- 1350
		x"00", -- 1351
		x"00", -- 1352
		x"00", -- 1353
		x"00", -- 1354
		x"00", -- 1355
		x"00", -- 1356
		x"00", -- 1357
		x"00", -- 1358
		x"00", -- 1359
		x"00", -- 135a
		x"30", -- 135b
		x"30", -- 135c
		x"10", -- 135d
		x"20", -- 135e
		x"00", -- 135f
		x"00", -- 1360
		x"00", -- 1361
		x"00", -- 1362
		x"00", -- 1363
		x"00", -- 1364
		x"00", -- 1365
		x"00", -- 1366
		x"00", -- 1367
		x"30", -- 1368
		x"30", -- 1369
		x"00", -- 136a
		x"00", -- 136b
		x"00", -- 136c
		x"00", -- 136d
		x"00", -- 136e
		x"00", -- 136f
		x"00", -- 1370
		x"00", -- 1371
		x"00", -- 1372
		x"00", -- 1373
		x"00", -- 1374
		x"7f", -- 1375
		x"01", -- 1376
		x"01", -- 1377
		x"7f", -- 1378
		x"01", -- 1379
		x"02", -- 137a
		x"04", -- 137b
		x"18", -- 137c
		x"00", -- 137d
		x"00", -- 137e
		x"00", -- 137f
		x"00", -- 1380
		x"00", -- 1381
		x"00", -- 1382
		x"00", -- 1383
		x"00", -- 1384
		x"00", -- 1385
		x"00", -- 1386
		x"7c", -- 1387
		x"04", -- 1388
		x"18", -- 1389
		x"10", -- 138a
		x"10", -- 138b
		x"20", -- 138c
		x"00", -- 138d
		x"00", -- 138e
		x"00", -- 138f
		x"00", -- 1390
		x"00", -- 1391
		x"00", -- 1392
		x"00", -- 1393
		x"00", -- 1394
		x"00", -- 1395
		x"00", -- 1396
		x"04", -- 1397
		x"08", -- 1398
		x"18", -- 1399
		x"28", -- 139a
		x"08", -- 139b
		x"08", -- 139c
		x"00", -- 139d
		x"00", -- 139e
		x"00", -- 139f
		x"00", -- 13a0
		x"00", -- 13a1
		x"00", -- 13a2
		x"00", -- 13a3
		x"00", -- 13a4
		x"00", -- 13a5
		x"00", -- 13a6
		x"10", -- 13a7
		x"7c", -- 13a8
		x"44", -- 13a9
		x"04", -- 13aa
		x"08", -- 13ab
		x"10", -- 13ac
		x"00", -- 13ad
		x"00", -- 13ae
		x"00", -- 13af
		x"00", -- 13b0
		x"00", -- 13b1
		x"00", -- 13b2
		x"00", -- 13b3
		x"00", -- 13b4
		x"00", -- 13b5
		x"00", -- 13b6
		x"00", -- 13b7
		x"7c", -- 13b8
		x"10", -- 13b9
		x"10", -- 13ba
		x"10", -- 13bb
		x"7c", -- 13bc
		x"00", -- 13bd
		x"00", -- 13be
		x"00", -- 13bf
		x"00", -- 13c0
		x"00", -- 13c1
		x"00", -- 13c2
		x"00", -- 13c3
		x"00", -- 13c4
		x"00", -- 13c5
		x"00", -- 13c6
		x"08", -- 13c7
		x"7c", -- 13c8
		x"08", -- 13c9
		x"18", -- 13ca
		x"28", -- 13cb
		x"48", -- 13cc
		x"00", -- 13cd
		x"00", -- 13ce
		x"00", -- 13cf
		x"00", -- 13d0
		x"00", -- 13d1
		x"00", -- 13d2
		x"00", -- 13d3
		x"00", -- 13d4
		x"00", -- 13d5
		x"00", -- 13d6
		x"20", -- 13d7
		x"7c", -- 13d8
		x"24", -- 13d9
		x"28", -- 13da
		x"20", -- 13db
		x"20", -- 13dc
		x"00", -- 13dd
		x"00", -- 13de
		x"00", -- 13df
		x"00", -- 13e0
		x"00", -- 13e1
		x"00", -- 13e2
		x"00", -- 13e3
		x"00", -- 13e4
		x"00", -- 13e5
		x"00", -- 13e6
		x"00", -- 13e7
		x"38", -- 13e8
		x"08", -- 13e9
		x"08", -- 13ea
		x"08", -- 13eb
		x"7e", -- 13ec
		x"00", -- 13ed
		x"00", -- 13ee
		x"00", -- 13ef
		x"00", -- 13f0
		x"00", -- 13f1
		x"00", -- 13f2
		x"00", -- 13f3
		x"00", -- 13f4
		x"00", -- 13f5
		x"00", -- 13f6
		x"00", -- 13f7
		x"7c", -- 13f8
		x"04", -- 13f9
		x"3c", -- 13fa
		x"04", -- 13fb
		x"7c", -- 13fc
		x"00", -- 13fd
		x"00", -- 13fe
		x"00", -- 13ff
		x"00", -- 1400
		x"00", -- 1401
		x"00", -- 1402
		x"00", -- 1403
		x"00", -- 1404
		x"00", -- 1405
		x"00", -- 1406
		x"00", -- 1407
		x"54", -- 1408
		x"54", -- 1409
		x"04", -- 140a
		x"08", -- 140b
		x"10", -- 140c
		x"00", -- 140d
		x"00", -- 140e
		x"00", -- 140f
		x"00", -- 1410
		x"00", -- 1411
		x"00", -- 1412
		x"00", -- 1413
		x"00", -- 1414
		x"00", -- 1415
		x"00", -- 1416
		x"00", -- 1417
		x"7f", -- 1418
		x"00", -- 1419
		x"00", -- 141a
		x"00", -- 141b
		x"00", -- 141c
		x"00", -- 141d
		x"00", -- 141e
		x"00", -- 141f
		x"00", -- 1420
		x"00", -- 1421
		x"00", -- 1422
		x"00", -- 1423
		x"00", -- 1424
		x"7f", -- 1425
		x"01", -- 1426
		x"09", -- 1427
		x"0a", -- 1428
		x"0c", -- 1429
		x"08", -- 142a
		x"08", -- 142b
		x"10", -- 142c
		x"00", -- 142d
		x"00", -- 142e
		x"00", -- 142f
		x"00", -- 1430
		x"00", -- 1431
		x"00", -- 1432
		x"00", -- 1433
		x"02", -- 1434
		x"04", -- 1435
		x"08", -- 1436
		x"18", -- 1437
		x"28", -- 1438
		x"48", -- 1439
		x"08", -- 143a
		x"08", -- 143b
		x"08", -- 143c
		x"00", -- 143d
		x"00", -- 143e
		x"00", -- 143f
		x"00", -- 1440
		x"00", -- 1441
		x"00", -- 1442
		x"00", -- 1443
		x"08", -- 1444
		x"08", -- 1445
		x"7f", -- 1446
		x"41", -- 1447
		x"41", -- 1448
		x"01", -- 1449
		x"02", -- 144a
		x"04", -- 144b
		x"08", -- 144c
		x"00", -- 144d
		x"00", -- 144e
		x"00", -- 144f
		x"00", -- 1450
		x"00", -- 1451
		x"00", -- 1452
		x"00", -- 1453
		x"00", -- 1454
		x"3e", -- 1455
		x"08", -- 1456
		x"08", -- 1457
		x"08", -- 1458
		x"08", -- 1459
		x"08", -- 145a
		x"7f", -- 145b
		x"00", -- 145c
		x"00", -- 145d
		x"00", -- 145e
		x"00", -- 145f
		x"00", -- 1460
		x"00", -- 1461
		x"00", -- 1462
		x"00", -- 1463
		x"04", -- 1464
		x"04", -- 1465
		x"7f", -- 1466
		x"04", -- 1467
		x"0c", -- 1468
		x"14", -- 1469
		x"24", -- 146a
		x"44", -- 146b
		x"04", -- 146c
		x"00", -- 146d
		x"00", -- 146e
		x"00", -- 146f
		x"00", -- 1470
		x"00", -- 1471
		x"00", -- 1472
		x"00", -- 1473
		x"10", -- 1474
		x"10", -- 1475
		x"7f", -- 1476
		x"11", -- 1477
		x"11", -- 1478
		x"11", -- 1479
		x"11", -- 147a
		x"21", -- 147b
		x"42", -- 147c
		x"00", -- 147d
		x"00", -- 147e
		x"00", -- 147f
		x"00", -- 1480
		x"00", -- 1481
		x"00", -- 1482
		x"00", -- 1483
		x"08", -- 1484
		x"08", -- 1485
		x"3e", -- 1486
		x"08", -- 1487
		x"08", -- 1488
		x"7f", -- 1489
		x"08", -- 148a
		x"08", -- 148b
		x"08", -- 148c
		x"00", -- 148d
		x"00", -- 148e
		x"00", -- 148f
		x"00", -- 1490
		x"00", -- 1491
		x"00", -- 1492
		x"00", -- 1493
		x"00", -- 1494
		x"1f", -- 1495
		x"21", -- 1496
		x"41", -- 1497
		x"01", -- 1498
		x"02", -- 1499
		x"04", -- 149a
		x"08", -- 149b
		x"10", -- 149c
		x"00", -- 149d
		x"00", -- 149e
		x"00", -- 149f
		x"00", -- 14a0
		x"00", -- 14a1
		x"00", -- 14a2
		x"00", -- 14a3
		x"10", -- 14a4
		x"10", -- 14a5
		x"1f", -- 14a6
		x"24", -- 14a7
		x"44", -- 14a8
		x"04", -- 14a9
		x"04", -- 14aa
		x"08", -- 14ab
		x"10", -- 14ac
		x"00", -- 14ad
		x"00", -- 14ae
		x"00", -- 14af
		x"00", -- 14b0
		x"00", -- 14b1
		x"00", -- 14b2
		x"00", -- 14b3
		x"00", -- 14b4
		x"7c", -- 14b5
		x"02", -- 14b6
		x"02", -- 14b7
		x"02", -- 14b8
		x"02", -- 14b9
		x"02", -- 14ba
		x"7e", -- 14bb
		x"00", -- 14bc
		x"00", -- 14bd
		x"00", -- 14be
		x"00", -- 14bf
		x"00", -- 14c0
		x"00", -- 14c1
		x"00", -- 14c2
		x"00", -- 14c3
		x"22", -- 14c4
		x"22", -- 14c5
		x"7f", -- 14c6
		x"22", -- 14c7
		x"22", -- 14c8
		x"02", -- 14c9
		x"04", -- 14ca
		x"08", -- 14cb
		x"10", -- 14cc
		x"00", -- 14cd
		x"00", -- 14ce
		x"00", -- 14cf
		x"00", -- 14d0
		x"00", -- 14d1
		x"00", -- 14d2
		x"00", -- 14d3
		x"00", -- 14d4
		x"70", -- 14d5
		x"00", -- 14d6
		x"01", -- 14d7
		x"71", -- 14d8
		x"01", -- 14d9
		x"02", -- 14da
		x"04", -- 14db
		x"78", -- 14dc
		x"00", -- 14dd
		x"00", -- 14de
		x"00", -- 14df
		x"00", -- 14e0
		x"00", -- 14e1
		x"00", -- 14e2
		x"00", -- 14e3
		x"00", -- 14e4
		x"7f", -- 14e5
		x"01", -- 14e6
		x"02", -- 14e7
		x"04", -- 14e8
		x"08", -- 14e9
		x"14", -- 14ea
		x"22", -- 14eb
		x"41", -- 14ec
		x"00", -- 14ed
		x"00", -- 14ee
		x"00", -- 14ef
		x"00", -- 14f0
		x"00", -- 14f1
		x"00", -- 14f2
		x"00", -- 14f3
		x"20", -- 14f4
		x"20", -- 14f5
		x"7f", -- 14f6
		x"21", -- 14f7
		x"22", -- 14f8
		x"24", -- 14f9
		x"20", -- 14fa
		x"20", -- 14fb
		x"1f", -- 14fc
		x"00", -- 14fd
		x"00", -- 14fe
		x"00", -- 14ff
		x"00", -- 1500
		x"00", -- 1501
		x"00", -- 1502
		x"00", -- 1503
		x"00", -- 1504
		x"41", -- 1505
		x"21", -- 1506
		x"11", -- 1507
		x"01", -- 1508
		x"02", -- 1509
		x"04", -- 150a
		x"08", -- 150b
		x"10", -- 150c
		x"00", -- 150d
		x"00", -- 150e
		x"00", -- 150f
		x"00", -- 1510
		x"00", -- 1511
		x"00", -- 1512
		x"00", -- 1513
		x"00", -- 1514
		x"1f", -- 1515
		x"11", -- 1516
		x"21", -- 1517
		x"51", -- 1518
		x"0a", -- 1519
		x"04", -- 151a
		x"08", -- 151b
		x"10", -- 151c
		x"00", -- 151d
		x"00", -- 151e
		x"00", -- 151f
		x"00", -- 1520
		x"00", -- 1521
		x"00", -- 1522
		x"00", -- 1523
		x"02", -- 1524
		x"3c", -- 1525
		x"08", -- 1526
		x"08", -- 1527
		x"7f", -- 1528
		x"08", -- 1529
		x"08", -- 152a
		x"10", -- 152b
		x"20", -- 152c
		x"00", -- 152d
		x"00", -- 152e
		x"00", -- 152f
		x"00", -- 1530
		x"00", -- 1531
		x"00", -- 1532
		x"00", -- 1533
		x"00", -- 1534
		x"49", -- 1535
		x"49", -- 1536
		x"49", -- 1537
		x"01", -- 1538
		x"01", -- 1539
		x"02", -- 153a
		x"04", -- 153b
		x"08", -- 153c
		x"00", -- 153d
		x"00", -- 153e
		x"00", -- 153f
		x"00", -- 1540
		x"00", -- 1541
		x"00", -- 1542
		x"00", -- 1543
		x"00", -- 1544
		x"3e", -- 1545
		x"00", -- 1546
		x"7f", -- 1547
		x"08", -- 1548
		x"08", -- 1549
		x"08", -- 154a
		x"10", -- 154b
		x"20", -- 154c
		x"00", -- 154d
		x"00", -- 154e
		x"00", -- 154f
		x"00", -- 1550
		x"00", -- 1551
		x"00", -- 1552
		x"00", -- 1553
		x"10", -- 1554
		x"10", -- 1555
		x"10", -- 1556
		x"18", -- 1557
		x"14", -- 1558
		x"12", -- 1559
		x"10", -- 155a
		x"10", -- 155b
		x"10", -- 155c
		x"00", -- 155d
		x"00", -- 155e
		x"00", -- 155f
		x"00", -- 1560
		x"00", -- 1561
		x"00", -- 1562
		x"00", -- 1563
		x"08", -- 1564
		x"08", -- 1565
		x"7f", -- 1566
		x"08", -- 1567
		x"08", -- 1568
		x"08", -- 1569
		x"08", -- 156a
		x"10", -- 156b
		x"20", -- 156c
		x"00", -- 156d
		x"00", -- 156e
		x"00", -- 156f
		x"00", -- 1570
		x"00", -- 1571
		x"00", -- 1572
		x"00", -- 1573
		x"00", -- 1574
		x"3e", -- 1575
		x"00", -- 1576
		x"00", -- 1577
		x"00", -- 1578
		x"00", -- 1579
		x"00", -- 157a
		x"7f", -- 157b
		x"00", -- 157c
		x"00", -- 157d
		x"00", -- 157e
		x"00", -- 157f
		x"00", -- 1580
		x"00", -- 1581
		x"00", -- 1582
		x"00", -- 1583
		x"00", -- 1584
		x"7f", -- 1585
		x"01", -- 1586
		x"02", -- 1587
		x"14", -- 1588
		x"08", -- 1589
		x"14", -- 158a
		x"22", -- 158b
		x"40", -- 158c
		x"00", -- 158d
		x"00", -- 158e
		x"00", -- 158f
		x"00", -- 1590
		x"00", -- 1591
		x"00", -- 1592
		x"00", -- 1593
		x"08", -- 1594
		x"7f", -- 1595
		x"02", -- 1596
		x"04", -- 1597
		x"0c", -- 1598
		x"1c", -- 1599
		x"2a", -- 159a
		x"49", -- 159b
		x"08", -- 159c
		x"00", -- 159d
		x"00", -- 159e
		x"00", -- 159f
		x"00", -- 15a0
		x"00", -- 15a1
		x"00", -- 15a2
		x"00", -- 15a3
		x"00", -- 15a4
		x"02", -- 15a5
		x"02", -- 15a6
		x"02", -- 15a7
		x"02", -- 15a8
		x"04", -- 15a9
		x"08", -- 15aa
		x"10", -- 15ab
		x"20", -- 15ac
		x"00", -- 15ad
		x"00", -- 15ae
		x"00", -- 15af
		x"00", -- 15b0
		x"00", -- 15b1
		x"00", -- 15b2
		x"00", -- 15b3
		x"00", -- 15b4
		x"04", -- 15b5
		x"22", -- 15b6
		x"21", -- 15b7
		x"21", -- 15b8
		x"21", -- 15b9
		x"21", -- 15ba
		x"21", -- 15bb
		x"41", -- 15bc
		x"00", -- 15bd
		x"00", -- 15be
		x"00", -- 15bf
		x"00", -- 15c0
		x"00", -- 15c1
		x"00", -- 15c2
		x"00", -- 15c3
		x"40", -- 15c4
		x"40", -- 15c5
		x"40", -- 15c6
		x"7e", -- 15c7
		x"40", -- 15c8
		x"40", -- 15c9
		x"40", -- 15ca
		x"40", -- 15cb
		x"3e", -- 15cc
		x"00", -- 15cd
		x"00", -- 15ce
		x"00", -- 15cf
		x"00", -- 15d0
		x"00", -- 15d1
		x"00", -- 15d2
		x"00", -- 15d3
		x"00", -- 15d4
		x"7f", -- 15d5
		x"01", -- 15d6
		x"01", -- 15d7
		x"01", -- 15d8
		x"02", -- 15d9
		x"04", -- 15da
		x"08", -- 15db
		x"30", -- 15dc
		x"00", -- 15dd
		x"00", -- 15de
		x"00", -- 15df
		x"00", -- 15e0
		x"00", -- 15e1
		x"00", -- 15e2
		x"00", -- 15e3
		x"00", -- 15e4
		x"10", -- 15e5
		x"28", -- 15e6
		x"44", -- 15e7
		x"02", -- 15e8
		x"01", -- 15e9
		x"01", -- 15ea
		x"01", -- 15eb
		x"01", -- 15ec
		x"00", -- 15ed
		x"00", -- 15ee
		x"00", -- 15ef
		x"00", -- 15f0
		x"00", -- 15f1
		x"00", -- 15f2
		x"00", -- 15f3
		x"08", -- 15f4
		x"08", -- 15f5
		x"7f", -- 15f6
		x"08", -- 15f7
		x"08", -- 15f8
		x"2a", -- 15f9
		x"29", -- 15fa
		x"49", -- 15fb
		x"08", -- 15fc
		x"00", -- 15fd
		x"00", -- 15fe
		x"00", -- 15ff
		x"00", -- 1600
		x"00", -- 1601
		x"00", -- 1602
		x"00", -- 1603
		x"00", -- 1604
		x"7f", -- 1605
		x"01", -- 1606
		x"01", -- 1607
		x"02", -- 1608
		x"14", -- 1609
		x"08", -- 160a
		x"04", -- 160b
		x"02", -- 160c
		x"00", -- 160d
		x"00", -- 160e
		x"00", -- 160f
		x"00", -- 1610
		x"00", -- 1611
		x"00", -- 1612
		x"00", -- 1613
		x"00", -- 1614
		x"3c", -- 1615
		x"02", -- 1616
		x"00", -- 1617
		x"3c", -- 1618
		x"00", -- 1619
		x"00", -- 161a
		x"7e", -- 161b
		x"01", -- 161c
		x"00", -- 161d
		x"00", -- 161e
		x"00", -- 161f
		x"00", -- 1620
		x"00", -- 1621
		x"00", -- 1622
		x"00", -- 1623
		x"00", -- 1624
		x"04", -- 1625
		x"08", -- 1626
		x"10", -- 1627
		x"20", -- 1628
		x"40", -- 1629
		x"41", -- 162a
		x"7f", -- 162b
		x"00", -- 162c
		x"00", -- 162d
		x"00", -- 162e
		x"00", -- 162f
		x"00", -- 1630
		x"00", -- 1631
		x"00", -- 1632
		x"00", -- 1633
		x"00", -- 1634
		x"01", -- 1635
		x"01", -- 1636
		x"22", -- 1637
		x"14", -- 1638
		x"08", -- 1639
		x"14", -- 163a
		x"22", -- 163b
		x"40", -- 163c
		x"00", -- 163d
		x"00", -- 163e
		x"00", -- 163f
		x"00", -- 1640
		x"00", -- 1641
		x"00", -- 1642
		x"00", -- 1643
		x"00", -- 1644
		x"7f", -- 1645
		x"10", -- 1646
		x"10", -- 1647
		x"7f", -- 1648
		x"10", -- 1649
		x"10", -- 164a
		x"10", -- 164b
		x"0f", -- 164c
		x"00", -- 164d
		x"00", -- 164e
		x"00", -- 164f
		x"00", -- 1650
		x"00", -- 1651
		x"00", -- 1652
		x"00", -- 1653
		x"10", -- 1654
		x"10", -- 1655
		x"7f", -- 1656
		x"11", -- 1657
		x"12", -- 1658
		x"14", -- 1659
		x"10", -- 165a
		x"10", -- 165b
		x"10", -- 165c
		x"00", -- 165d
		x"00", -- 165e
		x"00", -- 165f
		x"00", -- 1660
		x"00", -- 1661
		x"00", -- 1662
		x"00", -- 1663
		x"00", -- 1664
		x"3c", -- 1665
		x"04", -- 1666
		x"04", -- 1667
		x"04", -- 1668
		x"04", -- 1669
		x"04", -- 166a
		x"7f", -- 166b
		x"00", -- 166c
		x"00", -- 166d
		x"00", -- 166e
		x"00", -- 166f
		x"00", -- 1670
		x"00", -- 1671
		x"00", -- 1672
		x"00", -- 1673
		x"00", -- 1674
		x"7f", -- 1675
		x"01", -- 1676
		x"01", -- 1677
		x"3f", -- 1678
		x"01", -- 1679
		x"01", -- 167a
		x"7f", -- 167b
		x"00", -- 167c
		x"00", -- 167d
		x"00", -- 167e
		x"00", -- 167f
		x"00", -- 1680
		x"00", -- 1681
		x"00", -- 1682
		x"00", -- 1683
		x"00", -- 1684
		x"3e", -- 1685
		x"00", -- 1686
		x"7f", -- 1687
		x"01", -- 1688
		x"01", -- 1689
		x"02", -- 168a
		x"04", -- 168b
		x"18", -- 168c
		x"00", -- 168d
		x"00", -- 168e
		x"00", -- 168f
		x"00", -- 1690
		x"00", -- 1691
		x"00", -- 1692
		x"00", -- 1693
		x"00", -- 1694
		x"22", -- 1695
		x"22", -- 1696
		x"22", -- 1697
		x"22", -- 1698
		x"22", -- 1699
		x"02", -- 169a
		x"04", -- 169b
		x"08", -- 169c
		x"00", -- 169d
		x"00", -- 169e
		x"00", -- 169f
		x"00", -- 16a0
		x"00", -- 16a1
		x"00", -- 16a2
		x"00", -- 16a3
		x"00", -- 16a4
		x"28", -- 16a5
		x"28", -- 16a6
		x"28", -- 16a7
		x"28", -- 16a8
		x"29", -- 16a9
		x"29", -- 16aa
		x"2a", -- 16ab
		x"4c", -- 16ac
		x"00", -- 16ad
		x"00", -- 16ae
		x"00", -- 16af
		x"00", -- 16b0
		x"00", -- 16b1
		x"00", -- 16b2
		x"00", -- 16b3
		x"00", -- 16b4
		x"20", -- 16b5
		x"20", -- 16b6
		x"20", -- 16b7
		x"20", -- 16b8
		x"21", -- 16b9
		x"22", -- 16ba
		x"24", -- 16bb
		x"38", -- 16bc
		x"00", -- 16bd
		x"00", -- 16be
		x"00", -- 16bf
		x"00", -- 16c0
		x"00", -- 16c1
		x"00", -- 16c2
		x"00", -- 16c3
		x"00", -- 16c4
		x"3c", -- 16c5
		x"42", -- 16c6
		x"42", -- 16c7
		x"42", -- 16c8
		x"42", -- 16c9
		x"42", -- 16ca
		x"7e", -- 16cb
		x"00", -- 16cc
		x"00", -- 16cd
		x"00", -- 16ce
		x"00", -- 16cf
		x"00", -- 16d0
		x"00", -- 16d1
		x"00", -- 16d2
		x"00", -- 16d3
		x"00", -- 16d4
		x"7f", -- 16d5
		x"41", -- 16d6
		x"41", -- 16d7
		x"01", -- 16d8
		x"01", -- 16d9
		x"02", -- 16da
		x"04", -- 16db
		x"18", -- 16dc
		x"00", -- 16dd
		x"00", -- 16de
		x"00", -- 16df
		x"00", -- 16e0
		x"00", -- 16e1
		x"00", -- 16e2
		x"00", -- 16e3
		x"00", -- 16e4
		x"00", -- 16e5
		x"70", -- 16e6
		x"01", -- 16e7
		x"01", -- 16e8
		x"02", -- 16e9
		x"04", -- 16ea
		x"08", -- 16eb
		x"70", -- 16ec
		x"00", -- 16ed
		x"00", -- 16ee
		x"00", -- 16ef
		x"00", -- 16f0
		x"00", -- 16f1
		x"48", -- 16f2
		x"48", -- 16f3
		x"48", -- 16f4
		x"00", -- 16f5
		x"00", -- 16f6
		x"00", -- 16f7
		x"00", -- 16f8
		x"00", -- 16f9
		x"00", -- 16fa
		x"00", -- 16fb
		x"00", -- 16fc
		x"00", -- 16fd
		x"00", -- 16fe
		x"00", -- 16ff
		x"00", -- 1700
		x"00", -- 1701
		x"30", -- 1702
		x"48", -- 1703
		x"48", -- 1704
		x"30", -- 1705
		x"00", -- 1706
		x"00", -- 1707
		x"00", -- 1708
		x"00", -- 1709
		x"00", -- 170a
		x"00", -- 170b
		x"00", -- 170c
		x"00", -- 170d
		x"00", -- 170e
		x"00", -- 170f
		x"00", -- 1710
		x"00", -- 1711
		x"78", -- 1712
		x"40", -- 1713
		x"70", -- 1714
		x"40", -- 1715
		x"78", -- 1716
		x"00", -- 1717
		x"0c", -- 1718
		x"12", -- 1719
		x"12", -- 171a
		x"12", -- 171b
		x"0c", -- 171c
		x"00", -- 171d
		x"00", -- 171e
		x"00", -- 171f
		x"00", -- 1720
		x"00", -- 1721
		x"78", -- 1722
		x"40", -- 1723
		x"70", -- 1724
		x"40", -- 1725
		x"78", -- 1726
		x"00", -- 1727
		x"04", -- 1728
		x"0c", -- 1729
		x"04", -- 172a
		x"04", -- 172b
		x"0e", -- 172c
		x"00", -- 172d
		x"00", -- 172e
		x"00", -- 172f
		x"00", -- 1730
		x"00", -- 1731
		x"78", -- 1732
		x"40", -- 1733
		x"70", -- 1734
		x"40", -- 1735
		x"78", -- 1736
		x"00", -- 1737
		x"0c", -- 1738
		x"12", -- 1739
		x"04", -- 173a
		x"08", -- 173b
		x"1e", -- 173c
		x"00", -- 173d
		x"00", -- 173e
		x"00", -- 173f
		x"00", -- 1740
		x"00", -- 1741
		x"78", -- 1742
		x"40", -- 1743
		x"70", -- 1744
		x"40", -- 1745
		x"78", -- 1746
		x"00", -- 1747
		x"1c", -- 1748
		x"02", -- 1749
		x"0c", -- 174a
		x"02", -- 174b
		x"1c", -- 174c
		x"00", -- 174d
		x"00", -- 174e
		x"00", -- 174f
		x"00", -- 1750
		x"00", -- 1751
		x"78", -- 1752
		x"40", -- 1753
		x"70", -- 1754
		x"40", -- 1755
		x"78", -- 1756
		x"00", -- 1757
		x"14", -- 1758
		x"14", -- 1759
		x"1e", -- 175a
		x"04", -- 175b
		x"04", -- 175c
		x"00", -- 175d
		x"00", -- 175e
		x"00", -- 175f
		x"00", -- 1760
		x"00", -- 1761
		x"78", -- 1762
		x"40", -- 1763
		x"70", -- 1764
		x"40", -- 1765
		x"78", -- 1766
		x"00", -- 1767
		x"1e", -- 1768
		x"10", -- 1769
		x"1c", -- 176a
		x"02", -- 176b
		x"1c", -- 176c
		x"00", -- 176d
		x"00", -- 176e
		x"00", -- 176f
		x"00", -- 1770
		x"00", -- 1771
		x"78", -- 1772
		x"40", -- 1773
		x"70", -- 1774
		x"40", -- 1775
		x"78", -- 1776
		x"00", -- 1777
		x"0c", -- 1778
		x"10", -- 1779
		x"1c", -- 177a
		x"12", -- 177b
		x"0c", -- 177c
		x"00", -- 177d
		x"00", -- 177e
		x"00", -- 177f
		x"00", -- 1780
		x"00", -- 1781
		x"78", -- 1782
		x"40", -- 1783
		x"70", -- 1784
		x"40", -- 1785
		x"78", -- 1786
		x"00", -- 1787
		x"1e", -- 1788
		x"02", -- 1789
		x"04", -- 178a
		x"08", -- 178b
		x"10", -- 178c
		x"00", -- 178d
		x"00", -- 178e
		x"00", -- 178f
		x"00", -- 1790
		x"00", -- 1791
		x"78", -- 1792
		x"40", -- 1793
		x"70", -- 1794
		x"40", -- 1795
		x"78", -- 1796
		x"00", -- 1797
		x"0c", -- 1798
		x"12", -- 1799
		x"0c", -- 179a
		x"12", -- 179b
		x"0c", -- 179c
		x"00", -- 179d
		x"00", -- 179e
		x"00", -- 179f
		x"00", -- 17a0
		x"00", -- 17a1
		x"78", -- 17a2
		x"40", -- 17a3
		x"70", -- 17a4
		x"40", -- 17a5
		x"78", -- 17a6
		x"00", -- 17a7
		x"0c", -- 17a8
		x"12", -- 17a9
		x"0e", -- 17aa
		x"02", -- 17ab
		x"0c", -- 17ac
		x"00", -- 17ad
		x"00", -- 17ae
		x"00", -- 17af
		x"00", -- 17b0
		x"00", -- 17b1
		x"78", -- 17b2
		x"40", -- 17b3
		x"70", -- 17b4
		x"40", -- 17b5
		x"78", -- 17b6
		x"00", -- 17b7
		x"0c", -- 17b8
		x"12", -- 17b9
		x"1e", -- 17ba
		x"12", -- 17bb
		x"12", -- 17bc
		x"00", -- 17bd
		x"00", -- 17be
		x"00", -- 17bf
		x"00", -- 17c0
		x"00", -- 17c1
		x"78", -- 17c2
		x"40", -- 17c3
		x"70", -- 17c4
		x"40", -- 17c5
		x"78", -- 17c6
		x"00", -- 17c7
		x"1c", -- 17c8
		x"12", -- 17c9
		x"1c", -- 17ca
		x"12", -- 17cb
		x"1c", -- 17cc
		x"00", -- 17cd
		x"00", -- 17ce
		x"00", -- 17cf
		x"00", -- 17d0
		x"00", -- 17d1
		x"78", -- 17d2
		x"40", -- 17d3
		x"70", -- 17d4
		x"40", -- 17d5
		x"78", -- 17d6
		x"00", -- 17d7
		x"0e", -- 17d8
		x"10", -- 17d9
		x"10", -- 17da
		x"10", -- 17db
		x"0e", -- 17dc
		x"00", -- 17dd
		x"00", -- 17de
		x"00", -- 17df
		x"00", -- 17e0
		x"00", -- 17e1
		x"78", -- 17e2
		x"40", -- 17e3
		x"70", -- 17e4
		x"40", -- 17e5
		x"78", -- 17e6
		x"00", -- 17e7
		x"1c", -- 17e8
		x"12", -- 17e9
		x"12", -- 17ea
		x"12", -- 17eb
		x"1c", -- 17ec
		x"00", -- 17ed
		x"00", -- 17ee
		x"00", -- 17ef
		x"00", -- 17f0
		x"00", -- 17f1
		x"78", -- 17f2
		x"40", -- 17f3
		x"70", -- 17f4
		x"40", -- 17f5
		x"78", -- 17f6
		x"00", -- 17f7
		x"1e", -- 17f8
		x"10", -- 17f9
		x"1c", -- 17fa
		x"10", -- 17fb
		x"1e", -- 17fc
		x"00", -- 17fd
		x"00", -- 17fe
		x"00", -- 17ff
		x"00", -- 1800
		x"00", -- 1801
		x"78", -- 1802
		x"40", -- 1803
		x"70", -- 1804
		x"40", -- 1805
		x"78", -- 1806
		x"00", -- 1807
		x"1e", -- 1808
		x"10", -- 1809
		x"1c", -- 180a
		x"10", -- 180b
		x"10", -- 180c
		x"00", -- 180d
		x"00", -- 180e
		x"00", -- 180f
		x"00", -- 1810
		x"00", -- 1811
		x"78", -- 1812
		x"40", -- 1813
		x"70", -- 1814
		x"40", -- 1815
		x"40", -- 1816
		x"00", -- 1817
		x"0c", -- 1818
		x"12", -- 1819
		x"12", -- 181a
		x"12", -- 181b
		x"0c", -- 181c
		x"00", -- 181d
		x"00", -- 181e
		x"00", -- 181f
		x"00", -- 1820
		x"00", -- 1821
		x"78", -- 1822
		x"40", -- 1823
		x"70", -- 1824
		x"40", -- 1825
		x"40", -- 1826
		x"00", -- 1827
		x"04", -- 1828
		x"0c", -- 1829
		x"04", -- 182a
		x"04", -- 182b
		x"0e", -- 182c
		x"00", -- 182d
		x"00", -- 182e
		x"00", -- 182f
		x"00", -- 1830
		x"00", -- 1831
		x"78", -- 1832
		x"40", -- 1833
		x"70", -- 1834
		x"40", -- 1835
		x"40", -- 1836
		x"00", -- 1837
		x"0c", -- 1838
		x"12", -- 1839
		x"04", -- 183a
		x"08", -- 183b
		x"1e", -- 183c
		x"00", -- 183d
		x"00", -- 183e
		x"00", -- 183f
		x"00", -- 1840
		x"00", -- 1841
		x"78", -- 1842
		x"40", -- 1843
		x"70", -- 1844
		x"40", -- 1845
		x"40", -- 1846
		x"00", -- 1847
		x"1c", -- 1848
		x"02", -- 1849
		x"0c", -- 184a
		x"02", -- 184b
		x"1c", -- 184c
		x"00", -- 184d
		x"00", -- 184e
		x"00", -- 184f
		x"00", -- 1850
		x"00", -- 1851
		x"78", -- 1852
		x"40", -- 1853
		x"70", -- 1854
		x"40", -- 1855
		x"40", -- 1856
		x"00", -- 1857
		x"14", -- 1858
		x"14", -- 1859
		x"1e", -- 185a
		x"04", -- 185b
		x"04", -- 185c
		x"00", -- 185d
		x"00", -- 185e
		x"00", -- 185f
		x"00", -- 1860
		x"00", -- 1861
		x"70", -- 1862
		x"20", -- 1863
		x"20", -- 1864
		x"20", -- 1865
		x"70", -- 1866
		x"00", -- 1867
		x"0c", -- 1868
		x"12", -- 1869
		x"12", -- 186a
		x"12", -- 186b
		x"0c", -- 186c
		x"00", -- 186d
		x"00", -- 186e
		x"00", -- 186f
		x"00", -- 1870
		x"00", -- 1871
		x"78", -- 1872
		x"40", -- 1873
		x"70", -- 1874
		x"40", -- 1875
		x"40", -- 1876
		x"00", -- 1877
		x"0c", -- 1878
		x"10", -- 1879
		x"1c", -- 187a
		x"12", -- 187b
		x"0c", -- 187c
		x"00", -- 187d
		x"00", -- 187e
		x"00", -- 187f
		x"00", -- 1880
		x"00", -- 1881
		x"78", -- 1882
		x"40", -- 1883
		x"70", -- 1884
		x"40", -- 1885
		x"40", -- 1886
		x"00", -- 1887
		x"1e", -- 1888
		x"02", -- 1889
		x"04", -- 188a
		x"08", -- 188b
		x"10", -- 188c
		x"00", -- 188d
		x"00", -- 188e
		x"00", -- 188f
		x"00", -- 1890
		x"00", -- 1891
		x"78", -- 1892
		x"40", -- 1893
		x"70", -- 1894
		x"40", -- 1895
		x"40", -- 1896
		x"00", -- 1897
		x"0c", -- 1898
		x"12", -- 1899
		x"0c", -- 189a
		x"12", -- 189b
		x"0c", -- 189c
		x"00", -- 189d
		x"00", -- 189e
		x"00", -- 189f
		x"00", -- 18a0
		x"00", -- 18a1
		x"78", -- 18a2
		x"40", -- 18a3
		x"70", -- 18a4
		x"40", -- 18a5
		x"40", -- 18a6
		x"00", -- 18a7
		x"0c", -- 18a8
		x"12", -- 18a9
		x"0e", -- 18aa
		x"02", -- 18ab
		x"0c", -- 18ac
		x"00", -- 18ad
		x"00", -- 18ae
		x"00", -- 18af
		x"00", -- 18b0
		x"00", -- 18b1
		x"78", -- 18b2
		x"40", -- 18b3
		x"70", -- 18b4
		x"40", -- 18b5
		x"40", -- 18b6
		x"00", -- 18b7
		x"0c", -- 18b8
		x"12", -- 18b9
		x"1e", -- 18ba
		x"12", -- 18bb
		x"12", -- 18bc
		x"00", -- 18bd
		x"00", -- 18be
		x"00", -- 18bf
		x"00", -- 18c0
		x"00", -- 18c1
		x"78", -- 18c2
		x"40", -- 18c3
		x"70", -- 18c4
		x"40", -- 18c5
		x"40", -- 18c6
		x"00", -- 18c7
		x"1c", -- 18c8
		x"12", -- 18c9
		x"1c", -- 18ca
		x"12", -- 18cb
		x"1c", -- 18cc
		x"00", -- 18cd
		x"00", -- 18ce
		x"00", -- 18cf
		x"00", -- 18d0
		x"00", -- 18d1
		x"78", -- 18d2
		x"40", -- 18d3
		x"70", -- 18d4
		x"40", -- 18d5
		x"40", -- 18d6
		x"00", -- 18d7
		x"0e", -- 18d8
		x"10", -- 18d9
		x"10", -- 18da
		x"10", -- 18db
		x"0e", -- 18dc
		x"00", -- 18dd
		x"00", -- 18de
		x"00", -- 18df
		x"00", -- 18e0
		x"00", -- 18e1
		x"78", -- 18e2
		x"40", -- 18e3
		x"70", -- 18e4
		x"40", -- 18e5
		x"40", -- 18e6
		x"00", -- 18e7
		x"1c", -- 18e8
		x"12", -- 18e9
		x"12", -- 18ea
		x"12", -- 18eb
		x"1c", -- 18ec
		x"00", -- 18ed
		x"00", -- 18ee
		x"00", -- 18ef
		x"00", -- 18f0
		x"00", -- 18f1
		x"78", -- 18f2
		x"40", -- 18f3
		x"70", -- 18f4
		x"40", -- 18f5
		x"40", -- 18f6
		x"00", -- 18f7
		x"1e", -- 18f8
		x"10", -- 18f9
		x"1c", -- 18fa
		x"10", -- 18fb
		x"1e", -- 18fc
		x"00", -- 18fd
		x"00", -- 18fe
		x"00", -- 18ff
		x"00", -- 1900
		x"00", -- 1901
		x"00", -- 1902
		x"3c", -- 1903
		x"7e", -- 1904
		x"5a", -- 1905
		x"56", -- 1906
		x"4e", -- 1907
		x"4e", -- 1908
		x"56", -- 1909
		x"5a", -- 190a
		x"7e", -- 190b
		x"3c", -- 190c
		x"00", -- 190d
		x"00", -- 190e
		x"00", -- 190f
		x"00", -- 1910
		x"00", -- 1911
		x"00", -- 1912
		x"00", -- 1913
		x"00", -- 1914
		x"00", -- 1915
		x"00", -- 1916
		x"00", -- 1917
		x"00", -- 1918
		x"00", -- 1919
		x"00", -- 191a
		x"00", -- 191b
		x"00", -- 191c
		x"00", -- 191d
		x"00", -- 191e
		x"00", -- 191f
		x"00", -- 1920
		x"00", -- 1921
		x"00", -- 1922
		x"00", -- 1923
		x"00", -- 1924
		x"00", -- 1925
		x"00", -- 1926
		x"00", -- 1927
		x"00", -- 1928
		x"00", -- 1929
		x"00", -- 192a
		x"00", -- 192b
		x"00", -- 192c
		x"00", -- 192d
		x"00", -- 192e
		x"00", -- 192f
		x"00", -- 1930
		x"00", -- 1931
		x"00", -- 1932
		x"00", -- 1933
		x"00", -- 1934
		x"00", -- 1935
		x"00", -- 1936
		x"00", -- 1937
		x"00", -- 1938
		x"00", -- 1939
		x"00", -- 193a
		x"00", -- 193b
		x"00", -- 193c
		x"00", -- 193d
		x"00", -- 193e
		x"00", -- 193f
		x"00", -- 1940
		x"00", -- 1941
		x"00", -- 1942
		x"00", -- 1943
		x"00", -- 1944
		x"00", -- 1945
		x"00", -- 1946
		x"00", -- 1947
		x"00", -- 1948
		x"00", -- 1949
		x"00", -- 194a
		x"00", -- 194b
		x"00", -- 194c
		x"00", -- 194d
		x"00", -- 194e
		x"00", -- 194f
		x"00", -- 1950
		x"00", -- 1951
		x"00", -- 1952
		x"00", -- 1953
		x"00", -- 1954
		x"00", -- 1955
		x"00", -- 1956
		x"00", -- 1957
		x"00", -- 1958
		x"00", -- 1959
		x"00", -- 195a
		x"00", -- 195b
		x"00", -- 195c
		x"00", -- 195d
		x"00", -- 195e
		x"00", -- 195f
		x"00", -- 1960
		x"00", -- 1961
		x"00", -- 1962
		x"00", -- 1963
		x"00", -- 1964
		x"00", -- 1965
		x"00", -- 1966
		x"00", -- 1967
		x"00", -- 1968
		x"00", -- 1969
		x"00", -- 196a
		x"00", -- 196b
		x"00", -- 196c
		x"00", -- 196d
		x"00", -- 196e
		x"00", -- 196f
		x"00", -- 1970
		x"00", -- 1971
		x"00", -- 1972
		x"00", -- 1973
		x"00", -- 1974
		x"00", -- 1975
		x"00", -- 1976
		x"00", -- 1977
		x"00", -- 1978
		x"00", -- 1979
		x"00", -- 197a
		x"00", -- 197b
		x"00", -- 197c
		x"00", -- 197d
		x"00", -- 197e
		x"00", -- 197f
		x"00", -- 1980
		x"00", -- 1981
		x"00", -- 1982
		x"00", -- 1983
		x"00", -- 1984
		x"00", -- 1985
		x"00", -- 1986
		x"00", -- 1987
		x"00", -- 1988
		x"00", -- 1989
		x"00", -- 198a
		x"00", -- 198b
		x"00", -- 198c
		x"00", -- 198d
		x"00", -- 198e
		x"00", -- 198f
		x"00", -- 1990
		x"00", -- 1991
		x"00", -- 1992
		x"00", -- 1993
		x"00", -- 1994
		x"00", -- 1995
		x"00", -- 1996
		x"00", -- 1997
		x"00", -- 1998
		x"00", -- 1999
		x"00", -- 199a
		x"00", -- 199b
		x"00", -- 199c
		x"00", -- 199d
		x"00", -- 199e
		x"00", -- 199f
		x"00", -- 19a0
		x"00", -- 19a1
		x"00", -- 19a2
		x"00", -- 19a3
		x"00", -- 19a4
		x"00", -- 19a5
		x"00", -- 19a6
		x"00", -- 19a7
		x"00", -- 19a8
		x"00", -- 19a9
		x"00", -- 19aa
		x"00", -- 19ab
		x"00", -- 19ac
		x"00", -- 19ad
		x"00", -- 19ae
		x"00", -- 19af
		x"00", -- 19b0
		x"00", -- 19b1
		x"00", -- 19b2
		x"00", -- 19b3
		x"00", -- 19b4
		x"00", -- 19b5
		x"00", -- 19b6
		x"00", -- 19b7
		x"00", -- 19b8
		x"00", -- 19b9
		x"00", -- 19ba
		x"00", -- 19bb
		x"00", -- 19bc
		x"00", -- 19bd
		x"00", -- 19be
		x"00", -- 19bf
		x"00", -- 19c0
		x"00", -- 19c1
		x"00", -- 19c2
		x"00", -- 19c3
		x"00", -- 19c4
		x"00", -- 19c5
		x"00", -- 19c6
		x"00", -- 19c7
		x"00", -- 19c8
		x"00", -- 19c9
		x"00", -- 19ca
		x"00", -- 19cb
		x"00", -- 19cc
		x"00", -- 19cd
		x"00", -- 19ce
		x"00", -- 19cf
		x"00", -- 19d0
		x"00", -- 19d1
		x"00", -- 19d2
		x"00", -- 19d3
		x"00", -- 19d4
		x"00", -- 19d5
		x"00", -- 19d6
		x"00", -- 19d7
		x"00", -- 19d8
		x"00", -- 19d9
		x"00", -- 19da
		x"00", -- 19db
		x"00", -- 19dc
		x"00", -- 19dd
		x"00", -- 19de
		x"00", -- 19df
		x"00", -- 19e0
		x"00", -- 19e1
		x"00", -- 19e2
		x"00", -- 19e3
		x"00", -- 19e4
		x"00", -- 19e5
		x"00", -- 19e6
		x"00", -- 19e7
		x"00", -- 19e8
		x"00", -- 19e9
		x"00", -- 19ea
		x"00", -- 19eb
		x"00", -- 19ec
		x"00", -- 19ed
		x"00", -- 19ee
		x"00", -- 19ef
		x"00", -- 19f0
		x"00", -- 19f1
		x"00", -- 19f2
		x"00", -- 19f3
		x"00", -- 19f4
		x"00", -- 19f5
		x"00", -- 19f6
		x"00", -- 19f7
		x"00", -- 19f8
		x"00", -- 19f9
		x"00", -- 19fa
		x"00", -- 19fb
		x"00", -- 19fc
		x"00", -- 19fd
		x"00", -- 19fe
		x"00", -- 19ff
		x"00", -- 1a00
		x"00", -- 1a01
		x"00", -- 1a02
		x"00", -- 1a03
		x"00", -- 1a04
		x"00", -- 1a05
		x"00", -- 1a06
		x"00", -- 1a07
		x"00", -- 1a08
		x"00", -- 1a09
		x"00", -- 1a0a
		x"00", -- 1a0b
		x"00", -- 1a0c
		x"00", -- 1a0d
		x"00", -- 1a0e
		x"00", -- 1a0f
		x"00", -- 1a10
		x"00", -- 1a11
		x"00", -- 1a12
		x"00", -- 1a13
		x"00", -- 1a14
		x"00", -- 1a15
		x"00", -- 1a16
		x"00", -- 1a17
		x"00", -- 1a18
		x"00", -- 1a19
		x"00", -- 1a1a
		x"00", -- 1a1b
		x"00", -- 1a1c
		x"00", -- 1a1d
		x"00", -- 1a1e
		x"00", -- 1a1f
		x"00", -- 1a20
		x"00", -- 1a21
		x"00", -- 1a22
		x"00", -- 1a23
		x"00", -- 1a24
		x"00", -- 1a25
		x"00", -- 1a26
		x"00", -- 1a27
		x"00", -- 1a28
		x"00", -- 1a29
		x"00", -- 1a2a
		x"00", -- 1a2b
		x"00", -- 1a2c
		x"00", -- 1a2d
		x"00", -- 1a2e
		x"00", -- 1a2f
		x"00", -- 1a30
		x"00", -- 1a31
		x"00", -- 1a32
		x"00", -- 1a33
		x"00", -- 1a34
		x"00", -- 1a35
		x"00", -- 1a36
		x"00", -- 1a37
		x"00", -- 1a38
		x"00", -- 1a39
		x"00", -- 1a3a
		x"00", -- 1a3b
		x"00", -- 1a3c
		x"00", -- 1a3d
		x"00", -- 1a3e
		x"00", -- 1a3f
		x"00", -- 1a40
		x"00", -- 1a41
		x"00", -- 1a42
		x"00", -- 1a43
		x"00", -- 1a44
		x"00", -- 1a45
		x"00", -- 1a46
		x"00", -- 1a47
		x"00", -- 1a48
		x"00", -- 1a49
		x"00", -- 1a4a
		x"00", -- 1a4b
		x"00", -- 1a4c
		x"00", -- 1a4d
		x"00", -- 1a4e
		x"00", -- 1a4f
		x"00", -- 1a50
		x"00", -- 1a51
		x"00", -- 1a52
		x"00", -- 1a53
		x"00", -- 1a54
		x"00", -- 1a55
		x"00", -- 1a56
		x"00", -- 1a57
		x"00", -- 1a58
		x"00", -- 1a59
		x"00", -- 1a5a
		x"00", -- 1a5b
		x"00", -- 1a5c
		x"00", -- 1a5d
		x"00", -- 1a5e
		x"00", -- 1a5f
		x"00", -- 1a60
		x"00", -- 1a61
		x"00", -- 1a62
		x"00", -- 1a63
		x"00", -- 1a64
		x"00", -- 1a65
		x"00", -- 1a66
		x"00", -- 1a67
		x"00", -- 1a68
		x"00", -- 1a69
		x"00", -- 1a6a
		x"00", -- 1a6b
		x"00", -- 1a6c
		x"00", -- 1a6d
		x"00", -- 1a6e
		x"00", -- 1a6f
		x"00", -- 1a70
		x"00", -- 1a71
		x"00", -- 1a72
		x"00", -- 1a73
		x"00", -- 1a74
		x"00", -- 1a75
		x"00", -- 1a76
		x"00", -- 1a77
		x"00", -- 1a78
		x"00", -- 1a79
		x"00", -- 1a7a
		x"00", -- 1a7b
		x"00", -- 1a7c
		x"00", -- 1a7d
		x"00", -- 1a7e
		x"00", -- 1a7f
		x"00", -- 1a80
		x"00", -- 1a81
		x"00", -- 1a82
		x"00", -- 1a83
		x"00", -- 1a84
		x"00", -- 1a85
		x"00", -- 1a86
		x"00", -- 1a87
		x"00", -- 1a88
		x"00", -- 1a89
		x"00", -- 1a8a
		x"00", -- 1a8b
		x"00", -- 1a8c
		x"00", -- 1a8d
		x"00", -- 1a8e
		x"00", -- 1a8f
		x"00", -- 1a90
		x"00", -- 1a91
		x"00", -- 1a92
		x"00", -- 1a93
		x"00", -- 1a94
		x"00", -- 1a95
		x"00", -- 1a96
		x"00", -- 1a97
		x"00", -- 1a98
		x"00", -- 1a99
		x"00", -- 1a9a
		x"00", -- 1a9b
		x"00", -- 1a9c
		x"00", -- 1a9d
		x"00", -- 1a9e
		x"00", -- 1a9f
		x"00", -- 1aa0
		x"00", -- 1aa1
		x"00", -- 1aa2
		x"00", -- 1aa3
		x"00", -- 1aa4
		x"00", -- 1aa5
		x"00", -- 1aa6
		x"00", -- 1aa7
		x"00", -- 1aa8
		x"00", -- 1aa9
		x"00", -- 1aaa
		x"00", -- 1aab
		x"00", -- 1aac
		x"00", -- 1aad
		x"00", -- 1aae
		x"00", -- 1aaf
		x"00", -- 1ab0
		x"00", -- 1ab1
		x"00", -- 1ab2
		x"00", -- 1ab3
		x"00", -- 1ab4
		x"00", -- 1ab5
		x"00", -- 1ab6
		x"00", -- 1ab7
		x"00", -- 1ab8
		x"00", -- 1ab9
		x"00", -- 1aba
		x"00", -- 1abb
		x"00", -- 1abc
		x"00", -- 1abd
		x"00", -- 1abe
		x"00", -- 1abf
		x"00", -- 1ac0
		x"00", -- 1ac1
		x"00", -- 1ac2
		x"00", -- 1ac3
		x"00", -- 1ac4
		x"00", -- 1ac5
		x"00", -- 1ac6
		x"00", -- 1ac7
		x"00", -- 1ac8
		x"00", -- 1ac9
		x"00", -- 1aca
		x"00", -- 1acb
		x"00", -- 1acc
		x"00", -- 1acd
		x"00", -- 1ace
		x"00", -- 1acf
		x"00", -- 1ad0
		x"00", -- 1ad1
		x"00", -- 1ad2
		x"00", -- 1ad3
		x"00", -- 1ad4
		x"00", -- 1ad5
		x"00", -- 1ad6
		x"00", -- 1ad7
		x"00", -- 1ad8
		x"00", -- 1ad9
		x"00", -- 1ada
		x"00", -- 1adb
		x"00", -- 1adc
		x"00", -- 1add
		x"00", -- 1ade
		x"00", -- 1adf
		x"00", -- 1ae0
		x"00", -- 1ae1
		x"00", -- 1ae2
		x"00", -- 1ae3
		x"00", -- 1ae4
		x"00", -- 1ae5
		x"00", -- 1ae6
		x"00", -- 1ae7
		x"00", -- 1ae8
		x"00", -- 1ae9
		x"00", -- 1aea
		x"00", -- 1aeb
		x"00", -- 1aec
		x"00", -- 1aed
		x"00", -- 1aee
		x"00", -- 1aef
		x"00", -- 1af0
		x"00", -- 1af1
		x"00", -- 1af2
		x"00", -- 1af3
		x"00", -- 1af4
		x"00", -- 1af5
		x"00", -- 1af6
		x"00", -- 1af7
		x"00", -- 1af8
		x"00", -- 1af9
		x"00", -- 1afa
		x"00", -- 1afb
		x"00", -- 1afc
		x"00", -- 1afd
		x"00", -- 1afe
		x"00", -- 1aff
		x"00", -- 1b00
		x"00", -- 1b01
		x"00", -- 1b02
		x"00", -- 1b03
		x"00", -- 1b04
		x"00", -- 1b05
		x"00", -- 1b06
		x"00", -- 1b07
		x"00", -- 1b08
		x"00", -- 1b09
		x"00", -- 1b0a
		x"00", -- 1b0b
		x"00", -- 1b0c
		x"00", -- 1b0d
		x"00", -- 1b0e
		x"00", -- 1b0f
		x"00", -- 1b10
		x"00", -- 1b11
		x"00", -- 1b12
		x"00", -- 1b13
		x"00", -- 1b14
		x"00", -- 1b15
		x"00", -- 1b16
		x"00", -- 1b17
		x"00", -- 1b18
		x"00", -- 1b19
		x"00", -- 1b1a
		x"00", -- 1b1b
		x"00", -- 1b1c
		x"00", -- 1b1d
		x"00", -- 1b1e
		x"00", -- 1b1f
		x"00", -- 1b20
		x"00", -- 1b21
		x"00", -- 1b22
		x"00", -- 1b23
		x"00", -- 1b24
		x"00", -- 1b25
		x"00", -- 1b26
		x"00", -- 1b27
		x"00", -- 1b28
		x"00", -- 1b29
		x"00", -- 1b2a
		x"00", -- 1b2b
		x"00", -- 1b2c
		x"00", -- 1b2d
		x"00", -- 1b2e
		x"00", -- 1b2f
		x"00", -- 1b30
		x"00", -- 1b31
		x"00", -- 1b32
		x"00", -- 1b33
		x"00", -- 1b34
		x"00", -- 1b35
		x"00", -- 1b36
		x"00", -- 1b37
		x"00", -- 1b38
		x"00", -- 1b39
		x"00", -- 1b3a
		x"00", -- 1b3b
		x"00", -- 1b3c
		x"00", -- 1b3d
		x"00", -- 1b3e
		x"00", -- 1b3f
		x"00", -- 1b40
		x"00", -- 1b41
		x"00", -- 1b42
		x"00", -- 1b43
		x"00", -- 1b44
		x"00", -- 1b45
		x"00", -- 1b46
		x"00", -- 1b47
		x"00", -- 1b48
		x"00", -- 1b49
		x"00", -- 1b4a
		x"00", -- 1b4b
		x"00", -- 1b4c
		x"00", -- 1b4d
		x"00", -- 1b4e
		x"00", -- 1b4f
		x"00", -- 1b50
		x"00", -- 1b51
		x"00", -- 1b52
		x"00", -- 1b53
		x"00", -- 1b54
		x"00", -- 1b55
		x"00", -- 1b56
		x"00", -- 1b57
		x"00", -- 1b58
		x"00", -- 1b59
		x"00", -- 1b5a
		x"00", -- 1b5b
		x"00", -- 1b5c
		x"00", -- 1b5d
		x"00", -- 1b5e
		x"00", -- 1b5f
		x"00", -- 1b60
		x"00", -- 1b61
		x"00", -- 1b62
		x"00", -- 1b63
		x"00", -- 1b64
		x"00", -- 1b65
		x"00", -- 1b66
		x"00", -- 1b67
		x"00", -- 1b68
		x"00", -- 1b69
		x"00", -- 1b6a
		x"00", -- 1b6b
		x"00", -- 1b6c
		x"00", -- 1b6d
		x"00", -- 1b6e
		x"00", -- 1b6f
		x"00", -- 1b70
		x"00", -- 1b71
		x"00", -- 1b72
		x"00", -- 1b73
		x"00", -- 1b74
		x"00", -- 1b75
		x"00", -- 1b76
		x"00", -- 1b77
		x"00", -- 1b78
		x"00", -- 1b79
		x"00", -- 1b7a
		x"00", -- 1b7b
		x"00", -- 1b7c
		x"00", -- 1b7d
		x"00", -- 1b7e
		x"00", -- 1b7f
		x"00", -- 1b80
		x"00", -- 1b81
		x"00", -- 1b82
		x"00", -- 1b83
		x"00", -- 1b84
		x"00", -- 1b85
		x"00", -- 1b86
		x"00", -- 1b87
		x"00", -- 1b88
		x"00", -- 1b89
		x"00", -- 1b8a
		x"00", -- 1b8b
		x"00", -- 1b8c
		x"00", -- 1b8d
		x"00", -- 1b8e
		x"00", -- 1b8f
		x"00", -- 1b90
		x"00", -- 1b91
		x"00", -- 1b92
		x"00", -- 1b93
		x"00", -- 1b94
		x"00", -- 1b95
		x"00", -- 1b96
		x"00", -- 1b97
		x"00", -- 1b98
		x"00", -- 1b99
		x"00", -- 1b9a
		x"00", -- 1b9b
		x"00", -- 1b9c
		x"00", -- 1b9d
		x"00", -- 1b9e
		x"00", -- 1b9f
		x"00", -- 1ba0
		x"00", -- 1ba1
		x"00", -- 1ba2
		x"00", -- 1ba3
		x"00", -- 1ba4
		x"00", -- 1ba5
		x"00", -- 1ba6
		x"00", -- 1ba7
		x"00", -- 1ba8
		x"00", -- 1ba9
		x"00", -- 1baa
		x"00", -- 1bab
		x"00", -- 1bac
		x"00", -- 1bad
		x"00", -- 1bae
		x"00", -- 1baf
		x"00", -- 1bb0
		x"00", -- 1bb1
		x"00", -- 1bb2
		x"00", -- 1bb3
		x"00", -- 1bb4
		x"00", -- 1bb5
		x"00", -- 1bb6
		x"00", -- 1bb7
		x"00", -- 1bb8
		x"00", -- 1bb9
		x"00", -- 1bba
		x"00", -- 1bbb
		x"00", -- 1bbc
		x"00", -- 1bbd
		x"00", -- 1bbe
		x"00", -- 1bbf
		x"00", -- 1bc0
		x"00", -- 1bc1
		x"00", -- 1bc2
		x"00", -- 1bc3
		x"00", -- 1bc4
		x"00", -- 1bc5
		x"00", -- 1bc6
		x"00", -- 1bc7
		x"00", -- 1bc8
		x"00", -- 1bc9
		x"00", -- 1bca
		x"00", -- 1bcb
		x"00", -- 1bcc
		x"00", -- 1bcd
		x"00", -- 1bce
		x"00", -- 1bcf
		x"00", -- 1bd0
		x"00", -- 1bd1
		x"00", -- 1bd2
		x"00", -- 1bd3
		x"00", -- 1bd4
		x"00", -- 1bd5
		x"00", -- 1bd6
		x"00", -- 1bd7
		x"00", -- 1bd8
		x"00", -- 1bd9
		x"00", -- 1bda
		x"00", -- 1bdb
		x"00", -- 1bdc
		x"00", -- 1bdd
		x"00", -- 1bde
		x"00", -- 1bdf
		x"00", -- 1be0
		x"00", -- 1be1
		x"00", -- 1be2
		x"00", -- 1be3
		x"00", -- 1be4
		x"00", -- 1be5
		x"00", -- 1be6
		x"00", -- 1be7
		x"00", -- 1be8
		x"00", -- 1be9
		x"00", -- 1bea
		x"00", -- 1beb
		x"00", -- 1bec
		x"00", -- 1bed
		x"00", -- 1bee
		x"00", -- 1bef
		x"00", -- 1bf0
		x"00", -- 1bf1
		x"00", -- 1bf2
		x"00", -- 1bf3
		x"00", -- 1bf4
		x"00", -- 1bf5
		x"00", -- 1bf6
		x"00", -- 1bf7
		x"00", -- 1bf8
		x"00", -- 1bf9
		x"00", -- 1bfa
		x"00", -- 1bfb
		x"00", -- 1bfc
		x"00", -- 1bfd
		x"00", -- 1bfe
		x"00", -- 1bff
		x"00", -- 1c00
		x"00", -- 1c01
		x"00", -- 1c02
		x"00", -- 1c03
		x"00", -- 1c04
		x"00", -- 1c05
		x"00", -- 1c06
		x"00", -- 1c07
		x"00", -- 1c08
		x"00", -- 1c09
		x"00", -- 1c0a
		x"00", -- 1c0b
		x"00", -- 1c0c
		x"00", -- 1c0d
		x"00", -- 1c0e
		x"00", -- 1c0f
		x"00", -- 1c10
		x"00", -- 1c11
		x"00", -- 1c12
		x"00", -- 1c13
		x"00", -- 1c14
		x"00", -- 1c15
		x"00", -- 1c16
		x"00", -- 1c17
		x"00", -- 1c18
		x"00", -- 1c19
		x"00", -- 1c1a
		x"00", -- 1c1b
		x"00", -- 1c1c
		x"00", -- 1c1d
		x"00", -- 1c1e
		x"00", -- 1c1f
		x"00", -- 1c20
		x"00", -- 1c21
		x"00", -- 1c22
		x"00", -- 1c23
		x"00", -- 1c24
		x"00", -- 1c25
		x"00", -- 1c26
		x"00", -- 1c27
		x"00", -- 1c28
		x"00", -- 1c29
		x"00", -- 1c2a
		x"00", -- 1c2b
		x"00", -- 1c2c
		x"00", -- 1c2d
		x"00", -- 1c2e
		x"00", -- 1c2f
		x"00", -- 1c30
		x"00", -- 1c31
		x"00", -- 1c32
		x"00", -- 1c33
		x"00", -- 1c34
		x"00", -- 1c35
		x"00", -- 1c36
		x"00", -- 1c37
		x"00", -- 1c38
		x"00", -- 1c39
		x"00", -- 1c3a
		x"00", -- 1c3b
		x"00", -- 1c3c
		x"00", -- 1c3d
		x"00", -- 1c3e
		x"00", -- 1c3f
		x"00", -- 1c40
		x"00", -- 1c41
		x"00", -- 1c42
		x"00", -- 1c43
		x"00", -- 1c44
		x"00", -- 1c45
		x"00", -- 1c46
		x"00", -- 1c47
		x"00", -- 1c48
		x"00", -- 1c49
		x"00", -- 1c4a
		x"00", -- 1c4b
		x"00", -- 1c4c
		x"00", -- 1c4d
		x"00", -- 1c4e
		x"00", -- 1c4f
		x"00", -- 1c50
		x"00", -- 1c51
		x"00", -- 1c52
		x"00", -- 1c53
		x"00", -- 1c54
		x"00", -- 1c55
		x"00", -- 1c56
		x"00", -- 1c57
		x"00", -- 1c58
		x"00", -- 1c59
		x"00", -- 1c5a
		x"00", -- 1c5b
		x"00", -- 1c5c
		x"00", -- 1c5d
		x"00", -- 1c5e
		x"00", -- 1c5f
		x"00", -- 1c60
		x"00", -- 1c61
		x"00", -- 1c62
		x"00", -- 1c63
		x"00", -- 1c64
		x"00", -- 1c65
		x"00", -- 1c66
		x"00", -- 1c67
		x"00", -- 1c68
		x"00", -- 1c69
		x"00", -- 1c6a
		x"00", -- 1c6b
		x"00", -- 1c6c
		x"00", -- 1c6d
		x"00", -- 1c6e
		x"00", -- 1c6f
		x"00", -- 1c70
		x"00", -- 1c71
		x"00", -- 1c72
		x"00", -- 1c73
		x"00", -- 1c74
		x"00", -- 1c75
		x"00", -- 1c76
		x"00", -- 1c77
		x"00", -- 1c78
		x"00", -- 1c79
		x"00", -- 1c7a
		x"00", -- 1c7b
		x"00", -- 1c7c
		x"00", -- 1c7d
		x"00", -- 1c7e
		x"00", -- 1c7f
		x"00", -- 1c80
		x"00", -- 1c81
		x"00", -- 1c82
		x"00", -- 1c83
		x"00", -- 1c84
		x"00", -- 1c85
		x"00", -- 1c86
		x"00", -- 1c87
		x"00", -- 1c88
		x"00", -- 1c89
		x"00", -- 1c8a
		x"00", -- 1c8b
		x"00", -- 1c8c
		x"00", -- 1c8d
		x"00", -- 1c8e
		x"00", -- 1c8f
		x"00", -- 1c90
		x"00", -- 1c91
		x"00", -- 1c92
		x"00", -- 1c93
		x"00", -- 1c94
		x"00", -- 1c95
		x"00", -- 1c96
		x"00", -- 1c97
		x"00", -- 1c98
		x"00", -- 1c99
		x"00", -- 1c9a
		x"00", -- 1c9b
		x"00", -- 1c9c
		x"00", -- 1c9d
		x"00", -- 1c9e
		x"00", -- 1c9f
		x"00", -- 1ca0
		x"00", -- 1ca1
		x"00", -- 1ca2
		x"00", -- 1ca3
		x"00", -- 1ca4
		x"00", -- 1ca5
		x"00", -- 1ca6
		x"00", -- 1ca7
		x"00", -- 1ca8
		x"00", -- 1ca9
		x"00", -- 1caa
		x"00", -- 1cab
		x"00", -- 1cac
		x"00", -- 1cad
		x"00", -- 1cae
		x"00", -- 1caf
		x"00", -- 1cb0
		x"00", -- 1cb1
		x"00", -- 1cb2
		x"00", -- 1cb3
		x"00", -- 1cb4
		x"00", -- 1cb5
		x"00", -- 1cb6
		x"00", -- 1cb7
		x"00", -- 1cb8
		x"00", -- 1cb9
		x"00", -- 1cba
		x"00", -- 1cbb
		x"00", -- 1cbc
		x"00", -- 1cbd
		x"00", -- 1cbe
		x"00", -- 1cbf
		x"00", -- 1cc0
		x"00", -- 1cc1
		x"00", -- 1cc2
		x"00", -- 1cc3
		x"00", -- 1cc4
		x"00", -- 1cc5
		x"00", -- 1cc6
		x"00", -- 1cc7
		x"00", -- 1cc8
		x"00", -- 1cc9
		x"00", -- 1cca
		x"00", -- 1ccb
		x"00", -- 1ccc
		x"00", -- 1ccd
		x"00", -- 1cce
		x"00", -- 1ccf
		x"00", -- 1cd0
		x"00", -- 1cd1
		x"00", -- 1cd2
		x"00", -- 1cd3
		x"00", -- 1cd4
		x"00", -- 1cd5
		x"00", -- 1cd6
		x"00", -- 1cd7
		x"00", -- 1cd8
		x"00", -- 1cd9
		x"00", -- 1cda
		x"00", -- 1cdb
		x"00", -- 1cdc
		x"00", -- 1cdd
		x"00", -- 1cde
		x"00", -- 1cdf
		x"00", -- 1ce0
		x"00", -- 1ce1
		x"00", -- 1ce2
		x"00", -- 1ce3
		x"00", -- 1ce4
		x"00", -- 1ce5
		x"00", -- 1ce6
		x"00", -- 1ce7
		x"00", -- 1ce8
		x"00", -- 1ce9
		x"00", -- 1cea
		x"00", -- 1ceb
		x"00", -- 1cec
		x"00", -- 1ced
		x"00", -- 1cee
		x"00", -- 1cef
		x"00", -- 1cf0
		x"00", -- 1cf1
		x"00", -- 1cf2
		x"00", -- 1cf3
		x"00", -- 1cf4
		x"00", -- 1cf5
		x"00", -- 1cf6
		x"00", -- 1cf7
		x"00", -- 1cf8
		x"00", -- 1cf9
		x"00", -- 1cfa
		x"00", -- 1cfb
		x"00", -- 1cfc
		x"00", -- 1cfd
		x"00", -- 1cfe
		x"00", -- 1cff
		x"00", -- 1d00
		x"00", -- 1d01
		x"00", -- 1d02
		x"00", -- 1d03
		x"00", -- 1d04
		x"00", -- 1d05
		x"00", -- 1d06
		x"00", -- 1d07
		x"00", -- 1d08
		x"00", -- 1d09
		x"00", -- 1d0a
		x"00", -- 1d0b
		x"00", -- 1d0c
		x"00", -- 1d0d
		x"00", -- 1d0e
		x"00", -- 1d0f
		x"00", -- 1d10
		x"00", -- 1d11
		x"00", -- 1d12
		x"00", -- 1d13
		x"00", -- 1d14
		x"00", -- 1d15
		x"00", -- 1d16
		x"00", -- 1d17
		x"00", -- 1d18
		x"00", -- 1d19
		x"00", -- 1d1a
		x"00", -- 1d1b
		x"00", -- 1d1c
		x"00", -- 1d1d
		x"00", -- 1d1e
		x"00", -- 1d1f
		x"00", -- 1d20
		x"00", -- 1d21
		x"00", -- 1d22
		x"00", -- 1d23
		x"00", -- 1d24
		x"00", -- 1d25
		x"00", -- 1d26
		x"00", -- 1d27
		x"00", -- 1d28
		x"00", -- 1d29
		x"00", -- 1d2a
		x"00", -- 1d2b
		x"00", -- 1d2c
		x"00", -- 1d2d
		x"00", -- 1d2e
		x"00", -- 1d2f
		x"00", -- 1d30
		x"00", -- 1d31
		x"00", -- 1d32
		x"00", -- 1d33
		x"00", -- 1d34
		x"00", -- 1d35
		x"00", -- 1d36
		x"00", -- 1d37
		x"00", -- 1d38
		x"00", -- 1d39
		x"00", -- 1d3a
		x"00", -- 1d3b
		x"00", -- 1d3c
		x"00", -- 1d3d
		x"00", -- 1d3e
		x"00", -- 1d3f
		x"00", -- 1d40
		x"00", -- 1d41
		x"00", -- 1d42
		x"00", -- 1d43
		x"00", -- 1d44
		x"00", -- 1d45
		x"00", -- 1d46
		x"00", -- 1d47
		x"00", -- 1d48
		x"00", -- 1d49
		x"00", -- 1d4a
		x"00", -- 1d4b
		x"00", -- 1d4c
		x"00", -- 1d4d
		x"00", -- 1d4e
		x"00", -- 1d4f
		x"00", -- 1d50
		x"00", -- 1d51
		x"00", -- 1d52
		x"00", -- 1d53
		x"00", -- 1d54
		x"00", -- 1d55
		x"00", -- 1d56
		x"00", -- 1d57
		x"00", -- 1d58
		x"00", -- 1d59
		x"00", -- 1d5a
		x"00", -- 1d5b
		x"00", -- 1d5c
		x"00", -- 1d5d
		x"00", -- 1d5e
		x"00", -- 1d5f
		x"00", -- 1d60
		x"00", -- 1d61
		x"00", -- 1d62
		x"00", -- 1d63
		x"00", -- 1d64
		x"00", -- 1d65
		x"00", -- 1d66
		x"00", -- 1d67
		x"00", -- 1d68
		x"00", -- 1d69
		x"00", -- 1d6a
		x"00", -- 1d6b
		x"00", -- 1d6c
		x"00", -- 1d6d
		x"00", -- 1d6e
		x"00", -- 1d6f
		x"00", -- 1d70
		x"00", -- 1d71
		x"00", -- 1d72
		x"00", -- 1d73
		x"00", -- 1d74
		x"00", -- 1d75
		x"00", -- 1d76
		x"00", -- 1d77
		x"00", -- 1d78
		x"00", -- 1d79
		x"00", -- 1d7a
		x"00", -- 1d7b
		x"00", -- 1d7c
		x"00", -- 1d7d
		x"00", -- 1d7e
		x"00", -- 1d7f
		x"00", -- 1d80
		x"00", -- 1d81
		x"00", -- 1d82
		x"00", -- 1d83
		x"00", -- 1d84
		x"00", -- 1d85
		x"00", -- 1d86
		x"00", -- 1d87
		x"00", -- 1d88
		x"00", -- 1d89
		x"00", -- 1d8a
		x"00", -- 1d8b
		x"00", -- 1d8c
		x"00", -- 1d8d
		x"00", -- 1d8e
		x"00", -- 1d8f
		x"00", -- 1d90
		x"00", -- 1d91
		x"00", -- 1d92
		x"00", -- 1d93
		x"00", -- 1d94
		x"00", -- 1d95
		x"00", -- 1d96
		x"00", -- 1d97
		x"00", -- 1d98
		x"00", -- 1d99
		x"00", -- 1d9a
		x"00", -- 1d9b
		x"00", -- 1d9c
		x"00", -- 1d9d
		x"00", -- 1d9e
		x"00", -- 1d9f
		x"00", -- 1da0
		x"00", -- 1da1
		x"00", -- 1da2
		x"00", -- 1da3
		x"00", -- 1da4
		x"00", -- 1da5
		x"00", -- 1da6
		x"00", -- 1da7
		x"00", -- 1da8
		x"00", -- 1da9
		x"00", -- 1daa
		x"00", -- 1dab
		x"00", -- 1dac
		x"00", -- 1dad
		x"00", -- 1dae
		x"00", -- 1daf
		x"00", -- 1db0
		x"00", -- 1db1
		x"00", -- 1db2
		x"00", -- 1db3
		x"00", -- 1db4
		x"00", -- 1db5
		x"00", -- 1db6
		x"00", -- 1db7
		x"00", -- 1db8
		x"00", -- 1db9
		x"00", -- 1dba
		x"00", -- 1dbb
		x"00", -- 1dbc
		x"00", -- 1dbd
		x"00", -- 1dbe
		x"00", -- 1dbf
		x"00", -- 1dc0
		x"00", -- 1dc1
		x"00", -- 1dc2
		x"00", -- 1dc3
		x"00", -- 1dc4
		x"00", -- 1dc5
		x"00", -- 1dc6
		x"00", -- 1dc7
		x"00", -- 1dc8
		x"00", -- 1dc9
		x"00", -- 1dca
		x"00", -- 1dcb
		x"00", -- 1dcc
		x"00", -- 1dcd
		x"00", -- 1dce
		x"00", -- 1dcf
		x"00", -- 1dd0
		x"00", -- 1dd1
		x"00", -- 1dd2
		x"00", -- 1dd3
		x"00", -- 1dd4
		x"00", -- 1dd5
		x"00", -- 1dd6
		x"00", -- 1dd7
		x"00", -- 1dd8
		x"00", -- 1dd9
		x"00", -- 1dda
		x"00", -- 1ddb
		x"00", -- 1ddc
		x"00", -- 1ddd
		x"00", -- 1dde
		x"00", -- 1ddf
		x"00", -- 1de0
		x"00", -- 1de1
		x"00", -- 1de2
		x"00", -- 1de3
		x"00", -- 1de4
		x"00", -- 1de5
		x"00", -- 1de6
		x"00", -- 1de7
		x"00", -- 1de8
		x"00", -- 1de9
		x"00", -- 1dea
		x"00", -- 1deb
		x"00", -- 1dec
		x"00", -- 1ded
		x"00", -- 1dee
		x"00", -- 1def
		x"00", -- 1df0
		x"00", -- 1df1
		x"00", -- 1df2
		x"00", -- 1df3
		x"00", -- 1df4
		x"00", -- 1df5
		x"00", -- 1df6
		x"00", -- 1df7
		x"00", -- 1df8
		x"00", -- 1df9
		x"00", -- 1dfa
		x"00", -- 1dfb
		x"00", -- 1dfc
		x"00", -- 1dfd
		x"00", -- 1dfe
		x"00", -- 1dff
		x"00", -- 1e00
		x"00", -- 1e01
		x"00", -- 1e02
		x"00", -- 1e03
		x"00", -- 1e04
		x"00", -- 1e05
		x"00", -- 1e06
		x"00", -- 1e07
		x"00", -- 1e08
		x"00", -- 1e09
		x"00", -- 1e0a
		x"00", -- 1e0b
		x"00", -- 1e0c
		x"00", -- 1e0d
		x"00", -- 1e0e
		x"00", -- 1e0f
		x"00", -- 1e10
		x"00", -- 1e11
		x"00", -- 1e12
		x"00", -- 1e13
		x"00", -- 1e14
		x"00", -- 1e15
		x"00", -- 1e16
		x"00", -- 1e17
		x"00", -- 1e18
		x"00", -- 1e19
		x"00", -- 1e1a
		x"00", -- 1e1b
		x"00", -- 1e1c
		x"00", -- 1e1d
		x"00", -- 1e1e
		x"00", -- 1e1f
		x"00", -- 1e20
		x"00", -- 1e21
		x"00", -- 1e22
		x"00", -- 1e23
		x"00", -- 1e24
		x"00", -- 1e25
		x"00", -- 1e26
		x"00", -- 1e27
		x"00", -- 1e28
		x"00", -- 1e29
		x"00", -- 1e2a
		x"00", -- 1e2b
		x"00", -- 1e2c
		x"00", -- 1e2d
		x"00", -- 1e2e
		x"00", -- 1e2f
		x"00", -- 1e30
		x"00", -- 1e31
		x"00", -- 1e32
		x"00", -- 1e33
		x"00", -- 1e34
		x"00", -- 1e35
		x"00", -- 1e36
		x"00", -- 1e37
		x"00", -- 1e38
		x"00", -- 1e39
		x"00", -- 1e3a
		x"00", -- 1e3b
		x"00", -- 1e3c
		x"00", -- 1e3d
		x"00", -- 1e3e
		x"00", -- 1e3f
		x"00", -- 1e40
		x"00", -- 1e41
		x"00", -- 1e42
		x"00", -- 1e43
		x"00", -- 1e44
		x"00", -- 1e45
		x"00", -- 1e46
		x"00", -- 1e47
		x"00", -- 1e48
		x"00", -- 1e49
		x"00", -- 1e4a
		x"00", -- 1e4b
		x"00", -- 1e4c
		x"00", -- 1e4d
		x"00", -- 1e4e
		x"00", -- 1e4f
		x"00", -- 1e50
		x"00", -- 1e51
		x"00", -- 1e52
		x"00", -- 1e53
		x"00", -- 1e54
		x"00", -- 1e55
		x"00", -- 1e56
		x"00", -- 1e57
		x"00", -- 1e58
		x"00", -- 1e59
		x"00", -- 1e5a
		x"00", -- 1e5b
		x"00", -- 1e5c
		x"00", -- 1e5d
		x"00", -- 1e5e
		x"00", -- 1e5f
		x"00", -- 1e60
		x"00", -- 1e61
		x"00", -- 1e62
		x"00", -- 1e63
		x"00", -- 1e64
		x"00", -- 1e65
		x"00", -- 1e66
		x"00", -- 1e67
		x"00", -- 1e68
		x"00", -- 1e69
		x"00", -- 1e6a
		x"00", -- 1e6b
		x"00", -- 1e6c
		x"00", -- 1e6d
		x"00", -- 1e6e
		x"00", -- 1e6f
		x"00", -- 1e70
		x"00", -- 1e71
		x"00", -- 1e72
		x"00", -- 1e73
		x"00", -- 1e74
		x"00", -- 1e75
		x"00", -- 1e76
		x"00", -- 1e77
		x"00", -- 1e78
		x"00", -- 1e79
		x"00", -- 1e7a
		x"00", -- 1e7b
		x"00", -- 1e7c
		x"00", -- 1e7d
		x"00", -- 1e7e
		x"00", -- 1e7f
		x"00", -- 1e80
		x"00", -- 1e81
		x"00", -- 1e82
		x"00", -- 1e83
		x"00", -- 1e84
		x"00", -- 1e85
		x"00", -- 1e86
		x"00", -- 1e87
		x"00", -- 1e88
		x"00", -- 1e89
		x"00", -- 1e8a
		x"00", -- 1e8b
		x"00", -- 1e8c
		x"00", -- 1e8d
		x"00", -- 1e8e
		x"00", -- 1e8f
		x"00", -- 1e90
		x"00", -- 1e91
		x"00", -- 1e92
		x"00", -- 1e93
		x"00", -- 1e94
		x"00", -- 1e95
		x"00", -- 1e96
		x"00", -- 1e97
		x"00", -- 1e98
		x"00", -- 1e99
		x"00", -- 1e9a
		x"00", -- 1e9b
		x"00", -- 1e9c
		x"00", -- 1e9d
		x"00", -- 1e9e
		x"00", -- 1e9f
		x"00", -- 1ea0
		x"00", -- 1ea1
		x"00", -- 1ea2
		x"00", -- 1ea3
		x"00", -- 1ea4
		x"00", -- 1ea5
		x"00", -- 1ea6
		x"00", -- 1ea7
		x"00", -- 1ea8
		x"00", -- 1ea9
		x"00", -- 1eaa
		x"00", -- 1eab
		x"00", -- 1eac
		x"00", -- 1ead
		x"00", -- 1eae
		x"00", -- 1eaf
		x"00", -- 1eb0
		x"00", -- 1eb1
		x"00", -- 1eb2
		x"00", -- 1eb3
		x"00", -- 1eb4
		x"00", -- 1eb5
		x"00", -- 1eb6
		x"00", -- 1eb7
		x"00", -- 1eb8
		x"00", -- 1eb9
		x"00", -- 1eba
		x"00", -- 1ebb
		x"00", -- 1ebc
		x"00", -- 1ebd
		x"00", -- 1ebe
		x"00", -- 1ebf
		x"00", -- 1ec0
		x"00", -- 1ec1
		x"00", -- 1ec2
		x"00", -- 1ec3
		x"00", -- 1ec4
		x"00", -- 1ec5
		x"00", -- 1ec6
		x"00", -- 1ec7
		x"00", -- 1ec8
		x"00", -- 1ec9
		x"00", -- 1eca
		x"00", -- 1ecb
		x"00", -- 1ecc
		x"00", -- 1ecd
		x"00", -- 1ece
		x"00", -- 1ecf
		x"00", -- 1ed0
		x"00", -- 1ed1
		x"00", -- 1ed2
		x"00", -- 1ed3
		x"00", -- 1ed4
		x"00", -- 1ed5
		x"00", -- 1ed6
		x"00", -- 1ed7
		x"00", -- 1ed8
		x"00", -- 1ed9
		x"00", -- 1eda
		x"00", -- 1edb
		x"00", -- 1edc
		x"00", -- 1edd
		x"00", -- 1ede
		x"00", -- 1edf
		x"00", -- 1ee0
		x"00", -- 1ee1
		x"00", -- 1ee2
		x"00", -- 1ee3
		x"00", -- 1ee4
		x"00", -- 1ee5
		x"00", -- 1ee6
		x"00", -- 1ee7
		x"00", -- 1ee8
		x"00", -- 1ee9
		x"00", -- 1eea
		x"00", -- 1eeb
		x"00", -- 1eec
		x"00", -- 1eed
		x"00", -- 1eee
		x"00", -- 1eef
		x"00", -- 1ef0
		x"00", -- 1ef1
		x"00", -- 1ef2
		x"00", -- 1ef3
		x"00", -- 1ef4
		x"00", -- 1ef5
		x"00", -- 1ef6
		x"00", -- 1ef7
		x"00", -- 1ef8
		x"00", -- 1ef9
		x"00", -- 1efa
		x"00", -- 1efb
		x"00", -- 1efc
		x"00", -- 1efd
		x"00", -- 1efe
		x"00", -- 1eff
		x"00", -- 1f00
		x"00", -- 1f01
		x"00", -- 1f02
		x"00", -- 1f03
		x"00", -- 1f04
		x"00", -- 1f05
		x"00", -- 1f06
		x"00", -- 1f07
		x"00", -- 1f08
		x"00", -- 1f09
		x"00", -- 1f0a
		x"00", -- 1f0b
		x"00", -- 1f0c
		x"00", -- 1f0d
		x"00", -- 1f0e
		x"00", -- 1f0f
		x"00", -- 1f10
		x"00", -- 1f11
		x"00", -- 1f12
		x"00", -- 1f13
		x"00", -- 1f14
		x"00", -- 1f15
		x"00", -- 1f16
		x"00", -- 1f17
		x"00", -- 1f18
		x"00", -- 1f19
		x"00", -- 1f1a
		x"00", -- 1f1b
		x"00", -- 1f1c
		x"00", -- 1f1d
		x"00", -- 1f1e
		x"00", -- 1f1f
		x"00", -- 1f20
		x"00", -- 1f21
		x"00", -- 1f22
		x"00", -- 1f23
		x"00", -- 1f24
		x"00", -- 1f25
		x"00", -- 1f26
		x"00", -- 1f27
		x"00", -- 1f28
		x"00", -- 1f29
		x"00", -- 1f2a
		x"00", -- 1f2b
		x"00", -- 1f2c
		x"00", -- 1f2d
		x"00", -- 1f2e
		x"00", -- 1f2f
		x"00", -- 1f30
		x"00", -- 1f31
		x"00", -- 1f32
		x"00", -- 1f33
		x"00", -- 1f34
		x"00", -- 1f35
		x"00", -- 1f36
		x"00", -- 1f37
		x"00", -- 1f38
		x"00", -- 1f39
		x"00", -- 1f3a
		x"00", -- 1f3b
		x"00", -- 1f3c
		x"00", -- 1f3d
		x"00", -- 1f3e
		x"00", -- 1f3f
		x"00", -- 1f40
		x"00", -- 1f41
		x"00", -- 1f42
		x"00", -- 1f43
		x"00", -- 1f44
		x"00", -- 1f45
		x"00", -- 1f46
		x"00", -- 1f47
		x"00", -- 1f48
		x"00", -- 1f49
		x"00", -- 1f4a
		x"00", -- 1f4b
		x"00", -- 1f4c
		x"00", -- 1f4d
		x"00", -- 1f4e
		x"00", -- 1f4f
		x"00", -- 1f50
		x"00", -- 1f51
		x"00", -- 1f52
		x"00", -- 1f53
		x"00", -- 1f54
		x"00", -- 1f55
		x"00", -- 1f56
		x"00", -- 1f57
		x"00", -- 1f58
		x"00", -- 1f59
		x"00", -- 1f5a
		x"00", -- 1f5b
		x"00", -- 1f5c
		x"00", -- 1f5d
		x"00", -- 1f5e
		x"00", -- 1f5f
		x"00", -- 1f60
		x"00", -- 1f61
		x"00", -- 1f62
		x"00", -- 1f63
		x"00", -- 1f64
		x"00", -- 1f65
		x"00", -- 1f66
		x"00", -- 1f67
		x"00", -- 1f68
		x"00", -- 1f69
		x"00", -- 1f6a
		x"00", -- 1f6b
		x"00", -- 1f6c
		x"00", -- 1f6d
		x"00", -- 1f6e
		x"00", -- 1f6f
		x"00", -- 1f70
		x"00", -- 1f71
		x"00", -- 1f72
		x"00", -- 1f73
		x"00", -- 1f74
		x"00", -- 1f75
		x"00", -- 1f76
		x"00", -- 1f77
		x"00", -- 1f78
		x"00", -- 1f79
		x"00", -- 1f7a
		x"00", -- 1f7b
		x"00", -- 1f7c
		x"00", -- 1f7d
		x"00", -- 1f7e
		x"00", -- 1f7f
		x"00", -- 1f80
		x"00", -- 1f81
		x"00", -- 1f82
		x"00", -- 1f83
		x"00", -- 1f84
		x"00", -- 1f85
		x"00", -- 1f86
		x"00", -- 1f87
		x"00", -- 1f88
		x"00", -- 1f89
		x"00", -- 1f8a
		x"00", -- 1f8b
		x"00", -- 1f8c
		x"00", -- 1f8d
		x"00", -- 1f8e
		x"00", -- 1f8f
		x"00", -- 1f90
		x"00", -- 1f91
		x"00", -- 1f92
		x"00", -- 1f93
		x"00", -- 1f94
		x"00", -- 1f95
		x"00", -- 1f96
		x"00", -- 1f97
		x"00", -- 1f98
		x"00", -- 1f99
		x"00", -- 1f9a
		x"00", -- 1f9b
		x"00", -- 1f9c
		x"00", -- 1f9d
		x"00", -- 1f9e
		x"00", -- 1f9f
		x"00", -- 1fa0
		x"00", -- 1fa1
		x"00", -- 1fa2
		x"00", -- 1fa3
		x"00", -- 1fa4
		x"00", -- 1fa5
		x"00", -- 1fa6
		x"00", -- 1fa7
		x"00", -- 1fa8
		x"00", -- 1fa9
		x"00", -- 1faa
		x"00", -- 1fab
		x"00", -- 1fac
		x"00", -- 1fad
		x"00", -- 1fae
		x"00", -- 1faf
		x"00", -- 1fb0
		x"00", -- 1fb1
		x"00", -- 1fb2
		x"00", -- 1fb3
		x"00", -- 1fb4
		x"00", -- 1fb5
		x"00", -- 1fb6
		x"00", -- 1fb7
		x"00", -- 1fb8
		x"00", -- 1fb9
		x"00", -- 1fba
		x"00", -- 1fbb
		x"00", -- 1fbc
		x"00", -- 1fbd
		x"00", -- 1fbe
		x"00", -- 1fbf
		x"00", -- 1fc0
		x"00", -- 1fc1
		x"00", -- 1fc2
		x"00", -- 1fc3
		x"00", -- 1fc4
		x"00", -- 1fc5
		x"00", -- 1fc6
		x"00", -- 1fc7
		x"00", -- 1fc8
		x"00", -- 1fc9
		x"00", -- 1fca
		x"00", -- 1fcb
		x"00", -- 1fcc
		x"00", -- 1fcd
		x"00", -- 1fce
		x"00", -- 1fcf
		x"00", -- 1fd0
		x"00", -- 1fd1
		x"00", -- 1fd2
		x"00", -- 1fd3
		x"00", -- 1fd4
		x"00", -- 1fd5
		x"00", -- 1fd6
		x"00", -- 1fd7
		x"00", -- 1fd8
		x"00", -- 1fd9
		x"00", -- 1fda
		x"00", -- 1fdb
		x"00", -- 1fdc
		x"00", -- 1fdd
		x"00", -- 1fde
		x"00", -- 1fdf
		x"00", -- 1fe0
		x"00", -- 1fe1
		x"00", -- 1fe2
		x"00", -- 1fe3
		x"00", -- 1fe4
		x"00", -- 1fe5
		x"00", -- 1fe6
		x"00", -- 1fe7
		x"00", -- 1fe8
		x"00", -- 1fe9
		x"00", -- 1fea
		x"00", -- 1feb
		x"00", -- 1fec
		x"00", -- 1fed
		x"00", -- 1fee
		x"00", -- 1fef
		x"00", -- 1ff0
		x"00", -- 1ff1
		x"00", -- 1ff2
		x"00", -- 1ff3
		x"00", -- 1ff4
		x"00", -- 1ff5
		x"00", -- 1ff6
		x"00", -- 1ff7
		x"00", -- 1ff8
		x"00", -- 1ff9
		x"00", -- 1ffa
		x"00", -- 1ffb
		x"00", -- 1ffc
		x"00", -- 1ffd
		x"5b", -- 1ffe
		x"06"  -- 1fff
);

begin
romp: process(clk_i)
begin
	if (rising_edge(clk_i)) then
		data_o <= rom_i(to_integer(unsigned(addr_i)));
	end if;
end process;
end rtl;
