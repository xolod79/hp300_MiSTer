library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bootrom is
	generic(
		addr_width : integer := 32768;
		addr_bits  : integer := 15;
		data_width : integer := 32
        );
port(
    clk_i  : in std_logic;
    addr_i : in std_logic_vector(addr_bits-1 downto 0);
    data_o : out std_logic_vector(data_width-1 downto 0)
);
end bootrom;

architecture rtl of bootrom is

type rom_type is array (0 to addr_width-1) of std_logic_vector(data_width-1 downto 0);
signal rom_i : rom_type := (
		x"00000100", -- 0
		x"0000040c", -- 4
		x"00004bca", -- 8
		x"fffffff4", -- c
		x"ffffffee", -- 10
		x"ffffffe8", -- 14
		x"ffffffe2", -- 18
		x"ffffffdc", -- 1c
		x"ffffffd6", -- 20
		x"ffffffd0", -- 24
		x"ffffffca", -- 28
		x"ffffffc4", -- 2c
		x"fffffee6", -- 30
		x"fffffee6", -- 34
		x"fffffee6", -- 38
		x"fffffee6", -- 3c
		x"fffffee6", -- 40
		x"fffffee6", -- 44
		x"fffffee6", -- 48
		x"fffffee6", -- 4c
		x"fffffee6", -- 50
		x"fffffee6", -- 54
		x"fffffee6", -- 58
		x"fffffee6", -- 5c
		x"ffffff1c", -- 60
		x"ffffffbe", -- 64
		x"ffffffb8", -- 68
		x"ffffffb2", -- 6c
		x"ffffffac", -- 70
		x"ffffffa6", -- 74
		x"ffffffa0", -- 78
		x"ffffff9a", -- 7c
		x"ffffff94", -- 80
		x"ffffff8e", -- 84
		x"ffffff88", -- 88
		x"ffffff82", -- 8c
		x"ffffff7c", -- 90
		x"ffffff76", -- 94
		x"ffffff70", -- 98
		x"ffffff6a", -- 9c
		x"ffffff64", -- a0
		x"ffffff5e", -- a4
		x"ffffff58", -- a8
		x"ffffff52", -- ac
		x"ffffff4c", -- b0
		x"ffffff46", -- b4
		x"ffffff40", -- b8
		x"ffffff3a", -- bc
		x"fffffee0", -- c0
		x"fffffee0", -- c4
		x"fffffee0", -- c8
		x"fffffee0", -- cc
		x"fffffee0", -- d0
		x"fffffee0", -- d4
		x"fffffee0", -- d8
		x"fffffee6", -- dc
		x"fffffee6", -- e0
		x"fffffee6", -- e4
		x"fffffee6", -- e8
		x"fffffee6", -- ec
		x"fffffee6", -- f0
		x"fffffee6", -- f4
		x"fffffee6", -- f8
		x"fffffee6", -- fc
		x"ffffff16", -- 100
		x"ffffff10", -- 104
		x"ffffff0a", -- 108
		x"ffffff04", -- 10c
		x"fffffefe", -- 110
		x"fffffef8", -- 114
		x"fffffef2", -- 118
		x"fffffeec", -- 11c
		x"4efa785e", -- 120
		x"4efa784a", -- 124
		x"4efa783a", -- 128
		x"4efa7832", -- 12c
		x"4efa784e", -- 130
		x"4efa784a", -- 134
		x"4efa7846", -- 138
		x"4efa516a", -- 13c
		x"4efa427c", -- 140
		x"4efa7832", -- 144
		x"4efa53c6", -- 148
		x"4efa53a0", -- 14c
		x"4efa54f8", -- 150
		x"000065fc", -- 154
		x"4efa54f6", -- 158
		x"4efa62d4", -- 15c
		x"4efa62de", -- 160
		x"4efa62e8", -- 164
		x"4efa62f2", -- 168
		x"4efa62fc", -- 16c
		x"4efa471e", -- 170
		x"4efa471a", -- 174
		x"4efa471c", -- 178
		x"4efa4718", -- 17c
		x"4efa4714", -- 180
		x"4efa4710", -- 184
		x"4efa4c52", -- 188
		x"4efa4c56", -- 18c
		x"4efa4c5c", -- 190
		x"4efa4c64", -- 194
		x"4efa4c68", -- 198
		x"4efa0266", -- 19c
		x"4efa4a78", -- 1a0
		x"4efa3f1c", -- 1a4
		x"4efa48e0", -- 1a8
		x"4efa490c", -- 1ac
		x"00004d20", -- 1b0
		x"4efa4a26", -- 1b4
		x"4efa4bc0", -- 1b8
		x"4efa77ce", -- 1bc
		x"4efa3f34", -- 1c0
		x"4efa63aa", -- 1c4
		x"4efa66c2", -- 1c8
		x"4efa779a", -- 1cc
		x"4efa77a2", -- 1d0
		x"4efa7a3c", -- 1d4
		x"4efa7792", -- 1d8
		x"4efa777e", -- 1dc
		x"4efa7776", -- 1e0
		x"4efa7796", -- 1e4
		x"4efa77a0", -- 1e8
		x"00808000", -- 1ec
		x"00801d7c", -- 1f0
		x"fffff400", -- 1f4
		x"fffff406", -- 1f8
		x"fffff40c", -- 1fc
		x"fffff412", -- 200
		x"fffff418", -- 204
		x"fffff41e", -- 208
		x"fffff424", -- 20c
		x"fffff42a", -- 210
		x"fffff430", -- 214
		x"fffff436", -- 218
		x"fffff43c", -- 21c
		x"fffff442", -- 220
		x"fffff448", -- 224
		x"fffff44e", -- 228
		x"fffff454", -- 22c
		x"fffff45a", -- 230
		x"fffff460", -- 234
		x"fffff466", -- 238
		x"fffff46c", -- 23c
		x"fffff472", -- 240
		x"fffff478", -- 244
		x"fffff47e", -- 248
		x"fffff484", -- 24c
		x"fffff48a", -- 250
		x"fffff490", -- 254
		x"fffff496", -- 258
		x"fffff49c", -- 25c
		x"fffff4a2", -- 260
		x"fffff4a8", -- 264
		x"fffff4ae", -- 268
		x"fffff4b4", -- 26c
		x"fffff4ba", -- 270
		x"fffff4c0", -- 274
		x"fffff4c6", -- 278
		x"fffff4cc", -- 27c
		x"fffff4d2", -- 280
		x"fffff4d8", -- 284
		x"fffff4de", -- 288
		x"fffff4e4", -- 28c
		x"fffff4ea", -- 290
		x"fffff4f0", -- 294
		x"fffff4f6", -- 298
		x"fffff4fc", -- 29c
		x"fffff502", -- 2a0
		x"fffff508", -- 2a4
		x"fffff50e", -- 2a8
		x"fffff514", -- 2ac
		x"fffff51a", -- 2b0
		x"fffff520", -- 2b4
		x"fffff526", -- 2b8
		x"fffff52c", -- 2bc
		x"fffff532", -- 2c0
		x"fffff538", -- 2c4
		x"fffff53e", -- 2c8
		x"fffff544", -- 2cc
		x"fffff54a", -- 2d0
		x"fffff550", -- 2d4
		x"fffff556", -- 2d8
		x"fffff55c", -- 2dc
		x"fffff562", -- 2e0
		x"fffff568", -- 2e4
		x"fffff56e", -- 2e8
		x"fffff574", -- 2ec
		x"fffff57a", -- 2f0
		x"fffff580", -- 2f4
		x"fffff586", -- 2f8
		x"fffff58c", -- 2fc
		x"fffff592", -- 300
		x"fffff598", -- 304
		x"fffff59e", -- 308
		x"fffff5a4", -- 30c
		x"fffff5aa", -- 310
		x"fffff5b0", -- 314
		x"fffff5b6", -- 318
		x"fffff5bc", -- 31c
		x"fffff5c2", -- 320
		x"fffff5c8", -- 324
		x"fffff5ce", -- 328
		x"fffff5d4", -- 32c
		x"fffff5da", -- 330
		x"fffff5e0", -- 334
		x"fffff5e6", -- 338
		x"fffff5ec", -- 33c
		x"fffff5f2", -- 340
		x"fffff5f8", -- 344
		x"fffff5fe", -- 348
		x"fffff604", -- 34c
		x"fffff60a", -- 350
		x"fffff610", -- 354
		x"fffff616", -- 358
		x"fffff61c", -- 35c
		x"fffff622", -- 360
		x"fffff628", -- 364
		x"fffff62e", -- 368
		x"fffff634", -- 36c
		x"fffff63a", -- 370
		x"fffff640", -- 374
		x"fffff646", -- 378
		x"fffff64c", -- 37c
		x"fffff652", -- 380
		x"fffff658", -- 384
		x"fffff65e", -- 388
		x"fffff664", -- 38c
		x"fffff66a", -- 390
		x"fffff670", -- 394
		x"fffff676", -- 398
		x"fffff67c", -- 39c
		x"fffff682", -- 3a0
		x"fffff688", -- 3a4
		x"fffff68e", -- 3a8
		x"fffff694", -- 3ac
		x"fffff69a", -- 3b0
		x"fffff6a0", -- 3b4
		x"fffff6a6", -- 3b8
		x"fffff6ac", -- 3bc
		x"fffff6b2", -- 3c0
		x"fffff6b8", -- 3c4
		x"fffff6be", -- 3c8
		x"fffff6c4", -- 3cc
		x"fffff6ca", -- 3d0
		x"fffff6d0", -- 3d4
		x"fffff6d6", -- 3d8
		x"fffff6dc", -- 3dc
		x"fffff6e2", -- 3e0
		x"fffff6e8", -- 3e4
		x"fffff6ee", -- 3e8
		x"fffff6f4", -- 3ec
		x"fffff6fa", -- 3f0
		x"fffff700", -- 3f4
		x"fffff706", -- 3f8
		x"fffff70c", -- 3fc
		x"7a016056", -- 400
		x"7a026052", -- 404
		x"7a0d604e", -- 408
		x"4ff80000", -- 40c
		x"2c4f2a4e", -- 410
		x"284d264c", -- 414
		x"244b224a", -- 418
		x"20492008", -- 41c
		x"22002401", -- 420
		x"26022803", -- 424
		x"2a042c05", -- 428
		x"2e06be8f", -- 42c
		x"661abebc", -- 430
		x"aaaaaaaa", -- 434
		x"671e2e7c", -- 438
		x"55555555", -- 43c
		x"4a8767cc", -- 440
		x"2e7caaaa", -- 444
		x"aaaa60c4", -- 448
		x"13fc00fe", -- 44c
		x"0001ffff", -- 450
		x"4e722700", -- 454
		x"7a027c28", -- 458
		x"08850003", -- 45c
		x"671c2878", -- 460
		x"fed4082c", -- 464
		x"0001000b", -- 468
		x"670408c5", -- 46c
		x"0001082c", -- 470
		x"0000000a", -- 474
		x"670408c6", -- 478
		x"00104ff8", -- 47c
		x"0100287c", -- 480
		x"20000000", -- 484
		x"08c60011", -- 488
		x"4dfa0038", -- 48c
		x"203ceeee", -- 490
		x"11112200", -- 494
		x"24012602", -- 498
		x"28032e04", -- 49c
		x"2447264a", -- 4a0
		x"43f8c000", -- 4a4
		x"41f80000", -- 4a8
		x"48e0f930", -- 4ac
		x"b1c962f8", -- 4b0
		x"41f8ffff", -- 4b4
		x"203c0001", -- 4b8
		x"00004a10", -- 4bc
		x"91c0b1cc", -- 4c0
		x"62f84dfa", -- 4c4
		x"001c7e80", -- 4c8
		x"70ff13c7", -- 4cc
		x"0001ffff", -- 4d0
		x"26022403", -- 4d4
--		x"51c8fffa", -- 4d8
		x"4e714e71", -- 4d8 disable LED animation
		x"e207be00", -- 4dc
		x"66ece24f", -- 4e0
		x"08050000", -- 4e4
		x"662c4dfa", -- 4e8
		x"002a41f9", -- 4ec
		x"0051ffff", -- 4f0
		x"705a72a5", -- 4f4
		x"1080b010", -- 4f8
		x"66061081", -- 4fc
		x"b2106712", -- 500
		x"53883010", -- 504
		x"32005241", -- 508
		x"3081b050", -- 50c
		x"660408c6", -- 510
		x"00044dfa", -- 514
		x"00084a79", -- 518
		x"00500000", -- 51c
		x"4dfa0026", -- 520
		x"41f90047", -- 524
		x"800370c1", -- 528
		x"c0100c00", -- 52c
		x"00806614", -- 530
		x"70c110bc", -- 534
		x"007ec010", -- 538
		x"727f0c00", -- 53c
		x"00806604", -- 540
		x"08860005", -- 544
		x"08850002", -- 548
		x"670408c6", -- 54c
		x"00060885", -- 550
		x"00004dfa", -- 554
		x"00f20806", -- 558
		x"00046726", -- 55c
		x"41f90051", -- 560
		x"fffe3010", -- 564
		x"3200e049", -- 568
		x"827c0010", -- 56c
		x"c27c0017", -- 570
		x"8c010800", -- 574
		x"000f6600", -- 578
		x"009ae648", -- 57c
		x"c07c001f", -- 580
		x"60780806", -- 584
		x"0005662c", -- 588
		x"4dfa002a", -- 58c
		x"08390002", -- 590
		x"00478003", -- 594
		x"671e7004", -- 598
		x"08390000", -- 59c
		x"00478005", -- 5a0
		x"66025240", -- 5a4
		x"4dfa0054", -- 5a8
		x"4a390051", -- 5ac
		x"27048c3c", -- 5b0
		x"00046046", -- 5b4
		x"4dfa001e", -- 5b8
		x"52864240", -- 5bc
		x"4a390051", -- 5c0
		x"27047002", -- 5c4
		x"52860839", -- 5c8
		x"00070051", -- 5cc
		x"2704672a", -- 5d0
		x"52406026", -- 5d4
		x"4dfa0024", -- 5d8
		x"13fc000f", -- 5dc
		x"00510001", -- 5e0
		x"41f90051", -- 5e4
		x"0003725a", -- 5e8
		x"1081b210", -- 5ec
		x"660c72a5", -- 5f0
		x"1081b210", -- 5f4
		x"660408c5", -- 5f8
		x"00074dfa", -- 5fc
		x"004a0800", -- 600
		x"00006704", -- 604
		x"08c50000", -- 608
		x"424249fa", -- 60c
		x"00066000", -- 610
		x"4d22223c", -- 614
		x"00200020", -- 618
		x"41f90051", -- 61c
		x"a000343c", -- 620
		x"03ff20c1", -- 624
		x"51cafffc", -- 628
		x"4a790053", -- 62c
		x"80000806", -- 630
		x"00046712", -- 634
		x"7418c439", -- 638
		x"0051fffe", -- 63c
		x"670808b9", -- 640
		x"00000051", -- 644
		x"fffd1e3c", -- 648
		x"00fd4a47", -- 64c
		x"6b0613c7", -- 650
		x"0001ffff", -- 654
		x"43f80000", -- 658
		x"4bf8c000", -- 65c
		x"4dfa007a", -- 660
		x"74fe203c", -- 664
		x"eeee1111", -- 668
		x"223c8888", -- 66c
		x"77775242", -- 670
		x"c141e358", -- 674
		x"4840e358", -- 678
		x"48400802", -- 67c
		x"00016618", -- 680
		x"204949fa", -- 684
		x"ffeab2a0", -- 688
		x"60242080", -- 68c
-- disable upper RAM test (disabled)
		x"b1cd62f6", -- 690
--		x"b1cd4e71", -- 690
		x"0c401111", -- 694
		x"66d86036", -- 698
--		x"4e716036", -- 698
		x"204d49fa", -- 69c
		x"0002b290", -- 6a0
		x"600820c0", -- 6a4
		x"b1c966f6", -- 6a8
		x"60e667f6", -- 6ac
		x"600267da", -- 6b0
		x"26012810", -- 6b4
		x"bffc0000", -- 6b8
		x"01006208", -- 6bc
		x"530743fa", -- 6c0
		x"51e86022", -- 6c4
		x"58882a48", -- 6c8
		x"b3cd6702", -- 6cc
		x"4ed4bffc", -- 6d0
		x"00000100", -- 6d4
		x"633e4e75", -- 6d8
		x"bffc0000", -- 6dc
		x"010062e4", -- 6e0
		x"550743fa", -- 6e4
		x"51de4a47", -- 6e8
		x"6b0613c7", -- 6ec
		x"0001ffff", -- 6f0
		x"4dfa001e", -- 6f4
		x"41f90051", -- 6f8
		x"21a00806", -- 6fc
		x"00006706", -- 700
		x"41f90051", -- 704
		x"27044241", -- 708
		x"12196704", -- 70c
		x"30c160f8", -- 710
		x"4e722700", -- 714
		x"49f8f738", -- 718
		x"21ccfed4", -- 71c
		x"1945000b", -- 720
		x"4278fdc0", -- 724
		x"4238fed9", -- 728
		x"08ac0004", -- 72c
		x"000b11c6", -- 730
		x"fed24846", -- 734
		x"1946000a", -- 738
		x"2947009e", -- 73c
		x"422c00a1", -- 740
		x"4dfa0008", -- 744
		x"42390088", -- 748
		x"0000007c", -- 74c
		x"07000038", -- 750
		x"0008fed2", -- 754
		x"11fc00fa", -- 758
		x"feda51f8", -- 75c
		x"fdcd2878", -- 760
		x"fed408ec", -- 764
		x"0006000a", -- 768
		x"422c00a1", -- 76c
		x"4ff8fdac", -- 770
		x"6100446e", -- 774
		x"297c0000", -- 778
		x"0d7c0018", -- 77c
		x"297c0000", -- 780
		x"4020001c", -- 784
		x"297c0000", -- 788
		x"407c0020", -- 78c
		x"397c001c", -- 790
		x"0334297c", -- 794
		x"000000fc", -- 798
		x"002c297c", -- 79c
		x"00000140", -- 7a0
		x"001442ac", -- 7a4
		x"00104eb9", -- 7a8
		x"0000d4b8", -- 7ac
		x"70216100", -- 7b0
		x"46804eb9", -- 7b4
		x"0001891a", -- 7b8
		x"08380000", -- 7bc
		x"fed96704", -- 7c0
		x"6100468e", -- 7c4
		x"700541f9", -- 7c8
		x"00020000", -- 7cc
		x"43f90040", -- 7d0
		x"000045f8", -- 7d4
		x"40004dfa", -- 7d8
		x"004c2f08", -- 7dc
		x"2a4f0c50", -- 7e0
		x"f0ff6640", -- 7e4
		x"08280001", -- 7e8
		x"00036738", -- 7ec
		x"1028000c", -- 7f0
		x"743fc042", -- 7f4
		x"52401228", -- 7f8
		x"000dc242", -- 7fc
		x"b0016624", -- 800
		x"08280004", -- 804
		x"0003660e", -- 808
		x"28280012", -- 80c
		x"61004698", -- 810
		x"20574a40", -- 814
		x"660e7006", -- 818
		x"61004616", -- 81c
		x"d1e80004", -- 820
		x"4ea80004", -- 824
		x"2e4d205f", -- 828
		x"d1cab3c8", -- 82c
		x"66ac2878", -- 830
		x"fed47007", -- 834
		x"610045fa", -- 838
		x"4bec0018", -- 83c
		x"2a554a95", -- 840
		x"67122f0d", -- 844
		x"2a554e95", -- 848
		x"2a5f588d", -- 84c
		x"dbd56100", -- 850
		x"026860ea", -- 854
		x"2878fed4", -- 858
		x"082c0000", -- 85c
		x"005c6708", -- 860
		x"41fafba2", -- 864
		x"60003b54", -- 868
		x"4a78fdc0", -- 86c
		x"661243f8", -- 870
		x"fdc241fa", -- 874
		x"53fc6100", -- 878
		x"42704238", -- 87c
		x"fdcc6058", -- 880
		x"2878fed4", -- 884
		x"2978fdce", -- 888
		x"0010202c", -- 88c
		x"0014d1b8", -- 890
		x"fdce4e55", -- 894
		x"fff441ed", -- 898
		x"fff443f8", -- 89c
		x"fdc2700a", -- 8a0
		x"10c010d9", -- 8a4
		x"53406efa", -- 8a8
		x"0c200020", -- 8ac
		x"6608532d", -- 8b0
		x"fff467ac", -- 8b4
		x"60f208ec", -- 8b8
		x"0002000a", -- 8bc
		x"2f38fedc", -- 8c0
		x"486dfff4", -- 8c4
		x"61003834", -- 8c8
		x"41fa51fd", -- 8cc
		x"61004efa", -- 8d0
		x"4efafffe", -- 8d4
		x"00000000", -- 8d8
		x"2878fed4", -- 8dc
		x"41fa502c", -- 8e0
		x"61004ee6", -- 8e4
		x"08ac0006", -- 8e8
		x"000a6100", -- 8ec
		x"42042a6c", -- 8f0
		x"033006ac", -- 8f4
		x"fffffeda", -- 8f8
		x"0330487a", -- 8fc
		x"3a6a2b4f", -- 900
		x"fff642ac", -- 904
		x"033642ad", -- 908
		x"ffe670ff", -- 90c
		x"2b40fee0", -- 910
		x"50edfedc", -- 914
		x"21fce0ff", -- 918
		x"fffffedc", -- 91c
		x"422dffea", -- 920
		x"70ff2b40", -- 924
		x"fee0426d", -- 928
		x"fff4526d", -- 92c
		x"fff46d00", -- 930
		x"00d4266c", -- 934
		x"001c4a93", -- 938
		x"67f02f0b", -- 93c
		x"265350ed", -- 940
		x"ffe451ed", -- 944
		x"ffec6100", -- 948
		x"013e6100", -- 94c
		x"016c48e7", -- 950
		x"fff8554f", -- 954
		x"3f2dfff4", -- 958
		x"1f2dffe4", -- 95c
		x"486dfff0", -- 960
		x"486dffec", -- 964
		x"50e76100", -- 968
		x"658a4eab", -- 96c
		x"00006100", -- 970
		x"65964a1f", -- 974
		x"4cdf1fff", -- 978
		x"6700007e", -- 97c
		x"51edffe4", -- 980
		x"4a2dffea", -- 984
		x"66140cad", -- 988
		x"e0ffffff", -- 98c
		x"fff0670a", -- 990
		x"50edffea", -- 994
		x"21edfff0", -- 998
		x"fedc6100", -- 99c
		x"00ea6100", -- 9a0
		x"011843ed", -- 9a4
		x"fee441f8", -- 9a8
		x"fdc27004", -- 9ac
		x"12c06100", -- 9b0
		x"413848e7", -- 9b4
		x"fff8554f", -- 9b8
		x"486dfee4", -- 9bc
		x"61006534", -- 9c0
		x"4eab0004", -- 9c4
		x"61006540", -- 9c8
		x"4a1f4cdf", -- 9cc
		x"1fff6722", -- 9d0
		x"4a2dfee4", -- 9d4
		x"67126100", -- 9d8
		x"01224a2d", -- 9dc
		x"fee56708", -- 9e0
		x"082c0003", -- 9e4
		x"000b6706", -- 9e8
		x"61000332", -- 9ec
		x"67026124", -- 9f0
		x"60a8611a", -- 9f4
		x"6000ff50", -- 9f8
		x"6114265f", -- 9fc
		x"588bd7d3", -- a00
		x"6000ff34", -- a04
		x"3b7c0001", -- a08
		x"fff46000", -- a0c
		x"ff1e6100", -- a10
		x"030c670c", -- a14
		x"2f2dfff0", -- a18
		x"486dfee4", -- a1c
		x"6000fea6", -- a20
		x"4e75d27c", -- a24
		x"00303001", -- a28
		x"10c04e75", -- a2c
		x"48e7c000", -- a30
		x"42813200", -- a34
		x"82fc000a", -- a38
		x"66287020", -- a3c
		x"61ea4841", -- a40
		x"66247020", -- a44
		x"61e24cdf", -- a48
		x"00034e75", -- a4c
		x"48e7c000", -- a50
		x"42813200", -- a54
		x"82fc0064", -- a58
		x"671461c6", -- a5c
		x"484182fc", -- a60
		x"000a61be", -- a64
		x"484161ba", -- a68
		x"4cdf0003", -- a6c
		x"4e754841", -- a70
		x"82fc000a", -- a74
		x"67ee60ea", -- a78
		x"48e7c000", -- a7c
		x"42813200", -- a80
		x"82fc000a", -- a84
		x"60dc2f08", -- a88
		x"082c0002", -- a8c
		x"005c6724", -- a90
		x"4a2c00a9", -- a94
		x"670641fa", -- a98
		x"4ed86004", -- a9c
		x"41fa4eaf", -- aa0
		x"61004d26", -- aa4
		x"082c0002", -- aa8
		x"005c66f8", -- aac
		x"41fa4e5c", -- ab0
		x"61004d16", -- ab4
		x"205f4e75", -- ab8
		x"48e70008", -- abc
		x"2878fed4", -- ac0
		x"082c0005", -- ac4
		x"000a6706", -- ac8
		x"4eba4d1a", -- acc
		x"6008082c", -- ad0
		x"0007000a", -- ad4
		x"67044eba", -- ad8
		x"4d544cdf", -- adc
		x"10004e75", -- ae0
		x"225f201f", -- ae4
		x"52800880", -- ae8
		x"0000245f", -- aec
		x"2878fed4", -- af0
		x"91ac0330", -- af4
		x"24ac0330", -- af8
		x"4ed148e7", -- afc
		x"e0e04240", -- b00
		x"41edfee4", -- b04
		x"10105240", -- b08
		x"08000000", -- b0c
		x"67025240", -- b10
		x"226c0330", -- b14
		x"92c02949", -- b18
		x"033032d8", -- b1c
		x"55406efa", -- b20
		x"226c0330", -- b24
		x"92fc001e", -- b28
		x"29490330", -- b2c
		x"41ec0000", -- b30
		x"45e9000a", -- b34
		x"24d83490", -- b38
		x"41ec00ce", -- b3c
		x"45e90010", -- b40
		x"700634d8", -- b44
		x"51c8fffc", -- b48
		x"236dfff0", -- b4c
		x"00064a29", -- b50
		x"001f660c", -- b54
		x"42290005", -- b58
		x"42290004", -- b5c
		x"60000090", -- b60
		x"0ca9e0ff", -- b64
		x"ffff0006", -- b68
		x"66081369", -- b6c
		x"001f0005", -- b70
		x"602841fa", -- b74
		x"50f445e9", -- b78
		x"001f4241", -- b7c
		x"1229001e", -- b80
		x"4a416604", -- b84
		x"745a600e", -- b88
		x"141a5341", -- b8c
		x"10186706", -- b90
		x"b0026602", -- b94
		x"60ea1342", -- b98
		x"00051029", -- b9c
		x"00056b0c", -- ba0
		x"72c60300", -- ba4
		x"6706ea89", -- ba8
		x"01016606", -- bac
		x"137c005a", -- bb0
		x"00050ca9", -- bb4
		x"e0ffffff", -- bb8
		x"00066606", -- bbc
		x"42290004", -- bc0
		x"602c1229", -- bc4
		x"00054200", -- bc8
		x"206dffe6", -- bcc
		x"b0fc0000", -- bd0
		x"6716b228", -- bd4
		x"0005660a", -- bd8
		x"b0280004", -- bdc
		x"6c041028", -- be0
		x"00042068", -- be4
		x"000060e4", -- be8
		x"52401340", -- bec
		x"0004236d", -- bf0
		x"ffe60000", -- bf4
		x"2b49ffe6", -- bf8
		x"4aa90000", -- bfc
		x"66063b7c", -- c00
		x"0001feda", -- c04
		x"61282029", -- c08
		x"0006b0ad", -- c0c
		x"fee06714", -- c10
		x"2b40fee0", -- c14
		x"41f8fdd2", -- c18
		x"22006100", -- c1c
		x"57044218", -- c20
		x"6134610a", -- c24
		x"6100009c", -- c28
		x"4cdf0707", -- c2c
		x"4e75322d", -- c30
		x"feda302c", -- c34
		x"0046e248", -- c38
		x"52404eac", -- c3c
		x"003c526d", -- c40
		x"feda302c", -- c44
		x"00565540", -- c48
		x"b06dfeda", -- c4c
		x"6c063b7c", -- c50
		x"0001feda", -- c54
		x"4e7508ec", -- c58
		x"0006000a", -- c5c
		x"322c0046", -- c60
		x"e24941f8", -- c64
		x"fdd24240", -- c68
		x"1018670a", -- c6c
		x"53416d12", -- c70
		x"4eac0036", -- c74
		x"60f27020", -- c78
		x"53416d06", -- c7c
		x"4eac0036", -- c80
		x"60f6322d", -- c84
		x"feda0c41", -- c88
		x"00016606", -- c8c
		x"4a2dfedc", -- c90
		x"6624302c", -- c94
		x"0046e248", -- c98
		x"52404eac", -- c9c
		x"003c7020", -- ca0
		x"322c0046", -- ca4
		x"e2494eac", -- ca8
		x"00365341", -- cac
		x"6ef808ac", -- cb0
		x"0006000a", -- cb4
		x"4e7551ed", -- cb8
		x"fedc08ac", -- cbc
		x"0006000a", -- cc0
		x"4e7541f8", -- cc4
		x"fdd230fc", -- cc8
		x"20204a29", -- ccc
		x"00056720", -- cd0
		x"42401029", -- cd4
		x"00046100", -- cd8
		x"fd5410e9", -- cdc
		x"000510fc", -- ce0
		x"00200ca9", -- ce4
		x"e0ffffff", -- ce8
		x"00066604", -- cec
		x"72016010", -- cf0
		x"42411229", -- cf4
		x"001e0c41", -- cf8
		x"00f96f04", -- cfc
		x"323c00f9", -- d00
		x"45e9001f", -- d04
		x"4a126604", -- d08
		x"14bc0020", -- d0c
		x"4a416f06", -- d10
		x"10da5341", -- d14
		x"60f64218", -- d18
		x"6000ff3c", -- d1c
		x"342c032c", -- d20
		x"4a026750", -- d24
		x"206dffe6", -- d28
		x"b0fc0000", -- d2c
		x"6746b468", -- d30
		x"00046706", -- d34
		x"20680000", -- d38
		x"60ee45e8", -- d3c
		x"001e1028", -- d40
		x"001e5240", -- d44
		x"43edfee4", -- d48
		x"12da5340", -- d4c
		x"6efa2b68", -- d50
		x"0006fff0", -- d54
		x"45e8000a", -- d58
		x"43ec0000", -- d5c
		x"22da3292", -- d60
		x"45e80010", -- d64
		x"43ec00ce", -- d68
		x"700632da", -- d6c
		x"51c8fffc", -- d70
		x"50c04e75", -- d74
		x"51c04e75", -- d78
		x"00000e60", -- d7c
		x"00000004", -- d80
		x"00000eba", -- d84
		x"00000004", -- d88
		x"00000f48", -- d8c
		x"00000004", -- d90
		x"00000f90", -- d94
		x"00000004", -- d98
		x"0000100c", -- d9c
		x"00000004", -- da0
		x"00001026", -- da4
		x"00000004", -- da8
		x"00001070", -- dac
		x"00000004", -- db0
		x"0000508c", -- db4
		x"00000004", -- db8
		x"00001422", -- dbc
		x"00000004", -- dc0
		x"000014b6", -- dc4
		x"00000004", -- dc8
		x"00001808", -- dcc
		x"00000004", -- dd0
		x"00001760", -- dd4
		x"00000004", -- dd8
		x"00004a66", -- ddc
		x"00000004", -- de0
		x"000014f6", -- de4
		x"00000004", -- de8
		x"000193c0", -- dec
		x"00000004", -- df0
		x"000015e8", -- df4
		x"00000004", -- df8
		x"000015fc", -- dfc
		x"00000004", -- e00
		x"00001672", -- e04
		x"00000004", -- e08
		x"00004890", -- e0c
		x"00000004", -- e10
		x"0000175a", -- e14
		x"00000004", -- e18
		x"0000489c", -- e1c
		x"00000004", -- e20
		x"0000177a", -- e24
		x"00000004", -- e28
		x"00001de0", -- e2c
		x"00000004", -- e30
		x"00001ec2", -- e34
		x"00000004", -- e38
		x"00004e0a", -- e3c
		x"00000004", -- e40
		x"0000189e", -- e44
		x"00000004", -- e48
		x"00001cd2", -- e4c
		x"00000004", -- e50
		x"00003ed8", -- e54
		x"00000004", -- e58
		x"00000000", -- e5c
		x"4dfa000a", -- e60
		x"33fc0000", -- e64
		x"005f400e", -- e68
		x"4e750838", -- e6c
		x"0004feda", -- e70
		x"67182f00", -- e74
		x"0279ffdf", -- e78
		x"005f400e", -- e7c
		x"70004e7b", -- e80
		x"00024e7b", -- e84
		x"00024e71", -- e88
		x"201f4e75", -- e8c
		x"08380004", -- e90
		x"feda67f6", -- e94
		x"2f000079", -- e98
		x"0020005f", -- e9c
		x"400e7009", -- ea0
		x"60dc0838", -- ea4
		x"0004feda", -- ea8
		x"67e02f00", -- eac
		x"4e7a0002", -- eb0
		x"00000008", -- eb4
		x"60c808f8", -- eb8
		x"0002feda", -- ebc
		x"08b80004", -- ec0
		x"feda204f", -- ec4
		x"4267487a", -- ec8
		x"000640e7", -- ecc
		x"4e73bfc8", -- ed0
		x"2e48664e", -- ed4
		x"08b80002", -- ed8
		x"feda41f8", -- edc
		x"ffee2f20", -- ee0
		x"3f2030bc", -- ee4
		x"4ef9217c", -- ee8
		x"00000f28", -- eec
		x"00027000", -- ef0
		x"81c030df", -- ef4
		x"20dfb07c", -- ef8
		x"20146626", -- efc
		x"08f80004", -- f00
		x"feda4280", -- f04
		x"08c00009", -- f08
		x"4e7b0002", -- f0c
		x"4e7a1002", -- f10
		x"08010009", -- f14
		x"670c4280", -- f18
		x"4e7b0002", -- f1c
		x"08f80002", -- f20
		x"feda4e75", -- f24
		x"302f0006", -- f28
		x"4e734dfa", -- f2c
		x"00104a39", -- f30
		x"005f8003", -- f34
		x"08b80001", -- f38
		x"feda4e75", -- f3c
		x"08f80001", -- f40
		x"feda4e75", -- f44
		x"61e40838", -- f48
		x"0001feda", -- f4c
		x"663c41f9", -- f50
		x"005f8000", -- f54
		x"117c0000", -- f58
		x"0003117c", -- f5c
		x"00840001", -- f60
		x"117c0001", -- f64
		x"0003117c", -- f68
		x"00010001", -- f6c
		x"117c00ff", -- f70
		x"0009117c", -- f74
		x"00ff000b", -- f78
		x"117c00ff", -- f7c
		x"000d117c", -- f80
		x"00ff000f", -- f84
		x"117c0000", -- f88
		x"00014e75", -- f8c
		x"70206100", -- f90
		x"3ea00838", -- f94
		x"0001feda", -- f98
		x"6626203c", -- f9c
		x"00000014", -- fa0
		x"2f004857", -- fa4
		x"4eba4274", -- fa8
		x"48574eba", -- fac
		x"428e6b00", -- fb0
		x"001451c8", -- fb4
		x"fff44857", -- fb8
		x"4eba4280", -- fbc
		x"6b000006", -- fc0
		x"4e722700", -- fc4
		x"584f4e75", -- fc8
		x"2f00700e", -- fcc
		x"08380004", -- fd0
		x"feda671a", -- fd4
		x"102f000e", -- fd8
		x"e848103b", -- fdc
		x"001c2f97", -- fe0
		x"00002faf", -- fe4
		x"00040004", -- fe8
		x"dec0201f", -- fec
		x"4e750838", -- ff0
		x"0002feda", -- ff4
		x"67de60e6", -- ff8
		x"08080c00", -- ffc
		x"00000000", -- 1000
		x"3a14205c", -- 1004
		x"00000000", -- 1008
		x"4dfa0016", -- 100c
		x"0c794ef9", -- 1010
		x"00880000", -- 1014
		x"660a2878", -- 1018
		x"fed408ec", -- 101c
		x"0006000b", -- 1020
		x"4e757008", -- 1024
		x"61003e0a", -- 1028
		x"2a4f4dfa", -- 102c
		x"001e45f9", -- 1030
		x"00428003", -- 1034
		x"47f90042", -- 1038
		x"80017231", -- 103c
		x"700f6100", -- 1040
		x"54b46606", -- 1044
		x"700f6100", -- 1048
		x"54502e4d", -- 104c
		x"2878fed4", -- 1050
		x"082c0006", -- 1054
		x"000b6602", -- 1058
		x"4e70203c", -- 105c
		x"00000014", -- 1060
		x"4e7151c8", -- 1064
		x"fffc6100", -- 1068
		x"fede4e75", -- 106c
		x"70096100", -- 1070
		x"3dc02878", -- 1074
		x"fed44238", -- 1078
		x"fdcc08f8", -- 107c
		x"0007fdcc", -- 1080
		x"08b80007", -- 1084
		x"fed208ac", -- 1088
		x"0004005c", -- 108c
		x"08ac0005", -- 1090
		x"005c50ec", -- 1094
		x"00a6297c", -- 1098
		x"00800000", -- 109c
		x"00a242ac", -- 10a0
		x"0048207c", -- 10a4
		x"00560000", -- 10a8
		x"29480048", -- 10ac
		x"2a4f4dfa", -- 10b0
		x"01021028", -- 10b4
		x"0001c03c", -- 10b8
		x"001f0c00", -- 10bc
		x"00196600", -- 10c0
		x"00f20828", -- 10c4
		x"00060001", -- 10c8
		x"660000e8", -- 10cc
		x"4dfa006e", -- 10d0
		x"42800108", -- 10d4
		x"00854a80", -- 10d8
		x"67620838", -- 10dc
		x"0006fdcc", -- 10e0
		x"663c48e7", -- 10e4
		x"fffe082c", -- 10e8
		x"0004000b", -- 10ec
		x"661c224c", -- 10f0
		x"2a499bfc", -- 10f4
		x"00010800", -- 10f8
		x"700a6100", -- 10fc
		x"3d344eba", -- 1100
		x"3e8a4a00", -- 1104
		x"67046000", -- 1108
		x"3ae82878", -- 110c
		x"fed44eb9", -- 1110
		x"00007c5e", -- 1114
		x"08f80006", -- 1118
		x"fdcc4cdf", -- 111c
		x"7fff246c", -- 1120
		x"0048223c", -- 1124
		x"00000100", -- 1128
		x"700b6100", -- 112c
		x"3d044eb9", -- 1130
		x"00007ce2", -- 1134
		x"08380005", -- 1138
		x"fdcc6656", -- 113c
		x"4dfa0054", -- 1140
		x"2878fed4", -- 1144
		x"207c0056", -- 1148
		x"00002948", -- 114c
		x"0048702d", -- 1150
		x"61003cde", -- 1154
		x"61004daa", -- 1158
		x"082c0004", -- 115c
		x"005c6708", -- 1160
		x"702c6100", -- 1164
		x"3ccc602a", -- 1168
		x"700c6100", -- 116c
		x"3cc44dfa", -- 1170
		x"002208b8", -- 1174
		x"0007fdcc", -- 1178
		x"08f80007", -- 117c
		x"fed2283c", -- 1180
		x"00004000", -- 1184
		x"206c0048", -- 1188
		x"61003d4c", -- 118c
		x"4a436700", -- 1190
		x"016a6100", -- 1194
		x"3cbc2878", -- 1198
		x"fed408ec", -- 119c
		x"0004005c", -- 11a0
		x"08b80007", -- 11a4
		x"fed208f8", -- 11a8
		x"0007fdcc", -- 11ac
		x"42ac0048", -- 11b0
		x"2e4d2878", -- 11b4
		x"fed4082c", -- 11b8
		x"0001000a", -- 11bc
		x"6700013c", -- 11c0
		x"41f90100", -- 11c4
		x"0000323c", -- 11c8
		x"00842a4f", -- 11cc
		x"4dfa0114", -- 11d0
		x"10280001", -- 11d4
		x"c03c001f", -- 11d8
		x"0c000019", -- 11dc
		x"660000f0", -- 11e0
		x"08280006", -- 11e4
		x"00016600", -- 11e8
		x"00e6700d", -- 11ec
		x"61003c42", -- 11f0
		x"2878fed4", -- 11f4
		x"29480048", -- 11f8
		x"283c0000", -- 11fc
		x"4000102c", -- 1200
		x"005c48e7", -- 1204
		x"c0882a4f", -- 1208
		x"4dfa00ba", -- 120c
		x"22486100", -- 1210
		x"3cc64a43", -- 1214
		x"660000ae", -- 1218
		x"4dfa007a", -- 121c
		x"42800109", -- 1220
		x"00854a80", -- 1224
		x"676e4cdf", -- 1228
		x"11030838", -- 122c
		x"0006fdcc", -- 1230
		x"663c48e7", -- 1234
		x"fffe082c", -- 1238
		x"0004000b", -- 123c
		x"661c224c", -- 1240
		x"2a499bfc", -- 1244
		x"00010800", -- 1248
		x"700a6100", -- 124c
		x"3be44eba", -- 1250
		x"3d3a4a00", -- 1254
		x"67046000", -- 1258
		x"39982878", -- 125c
		x"fed44eb9", -- 1260
		x"00007c5e", -- 1264
		x"08f80006", -- 1268
		x"fdcc4cdf", -- 126c
		x"7fff700b", -- 1270
		x"61003bbe", -- 1274
		x"246c0048", -- 1278
		x"4eb90000", -- 127c
		x"7ce20838", -- 1280
		x"0005fdcc", -- 1284
		x"66482878", -- 1288
		x"fed4102c", -- 128c
		x"005c48e7", -- 1290
		x"c0882a4f", -- 1294
		x"08ac0004", -- 1298
		x"005c700d", -- 129c
		x"61003b92", -- 12a0
		x"4dfa0022", -- 12a4
		x"61004c5a", -- 12a8
		x"2878fed4", -- 12ac
		x"082c0004", -- 12b0
		x"005c6610", -- 12b4
		x"4cdf1103", -- 12b8
		x"1940005c", -- 12bc
		x"08b80007", -- 12c0
		x"fdcc6036", -- 12c4
		x"2e4d4cdf", -- 12c8
		x"11031940", -- 12cc
		x"005c4245", -- 12d0
		x"1a280101", -- 12d4
		x"e44d5245", -- 12d8
		x"d2457416", -- 12dc
		x"e5add1c5", -- 12e0
		x"600a2e4d", -- 12e4
		x"d1fc0040", -- 12e8
		x"00005241", -- 12ec
		x"b1fc2000", -- 12f0
		x"00006600", -- 12f4
		x"fed642ac", -- 12f8
		x"00484dfa", -- 12fc
		x"00b42a4f", -- 1300
		x"2878fed4", -- 1304
		x"08ac0005", -- 1308
		x"005c08ac", -- 130c
		x"0007005c", -- 1310
		x"702e6100", -- 1314
		x"3b1c43f9", -- 1318
		x"00510001", -- 131c
		x"12bc000c", -- 1320
		x"137c0000", -- 1324
		x"00024dfa", -- 1328
		x"f5ac7032", -- 132c
		x"610068e4", -- 1330
		x"4dfa007e", -- 1334
		x"45f90051", -- 1338
		x"a0011212", -- 133c
		x"76001412", -- 1340
		x"76ffb401", -- 1344
		x"666a43f9", -- 1348
		x"0051b001", -- 134c
		x"7eff6100", -- 1350
		x"3bb24a40", -- 1354
		x"66267006", -- 1358
		x"c038fed2", -- 135c
		x"72140101", -- 1360
		x"672445f9", -- 1364
		x"0051a002", -- 1368
		x"43f90051", -- 136c
		x"b0022e3c", -- 1370
		x"7f7f7f7f", -- 1374
		x"61003b8c", -- 1378
		x"4a40670a", -- 137c
		x"61003ad2", -- 1380
		x"08ec0005", -- 1384
		x"005c223c", -- 1388
		x"00200020", -- 138c
		x"41f90051", -- 1390
		x"a000343c", -- 1394
		x"03ff20c1", -- 1398
		x"51cafffc", -- 139c
		x"08380007", -- 13a0
		x"fdcc6722", -- 13a4
		x"61004ab8", -- 13a8
		x"08b80007", -- 13ac
		x"fdcc6016", -- 13b0
		x"2e4d08ec", -- 13b4
		x"0007005c", -- 13b8
		x"4aac0048", -- 13bc
		x"66086100", -- 13c0
		x"4e446100", -- 13c4
		x"63962878", -- 13c8
		x"fed4397c", -- 13cc
		x"0001032e", -- 13d0
		x"61005d7c", -- 13d4
		x"41fa45be", -- 13d8
		x"610043ee", -- 13dc
		x"48ec0018", -- 13e0
		x"00724dfa", -- 13e4
		x"00224a79", -- 13e8
		x"00538000", -- 13ec
		x"08380004", -- 13f0
		x"fed26712", -- 13f4
		x"7018c039", -- 13f8
		x"0051fffe", -- 13fc
		x"670808b9", -- 1400
		x"00000051", -- 1404
		x"fffd08b8", -- 1408
		x"0007fdcc", -- 140c
		x"0cac0000", -- 1410
		x"62080030", -- 1414
		x"660608f8", -- 1418
		x"0007fdcc", -- 141c
		x"4e75700e", -- 1420
		x"61003a0e", -- 1424
		x"41f80000", -- 1428
		x"283c0001", -- 142c
		x"c0004dfa", -- 1430
		x"001e224f", -- 1434
-- disable bootrom checksum
--		x"61003a70", -- 1438
		x"4e714e71", -- 1438
		x"082c0006", -- 143c
		x"000b6604", -- 1440
--		x"4a40660a", -- 1444
		x"4a40600a", -- 1444
		x"41fa2b86", -- 1448
		x"61003a32", -- 144c
		x"600a2e49", -- 1450
		x"41fa2b7a", -- 1454
		x"61003a2a", -- 1458
		x"2878fed4", -- 145c
		x"4cec0018", -- 1460
		x"0072702d", -- 1464
		x"610039ca", -- 1468
		x"082c0004", -- 146c
		x"005c670a", -- 1470
		x"41fa46c6", -- 1474
		x"61003a0a", -- 1478
		x"60100838", -- 147c
		x"0007fed2", -- 1480
		x"670841fa", -- 1484
		x"46b46100", -- 1488
		x"39f4702e", -- 148c
		x"610039a2", -- 1490
		x"41fa469a", -- 1494
		x"082c0007", -- 1498
		x"005c6614", -- 149c
		x"082c0005", -- 14a0
		x"005c6604", -- 14a4
		x"600039d6", -- 14a8
		x"610039d6", -- 14ac
		x"60003b6c", -- 14b0
		x"4e7541fa", -- 14b4
		x"466543f8", -- 14b8
		x"fdd212d8", -- 14bc
		x"66fc0838", -- 14c0
		x"0002feda", -- 14c4
		x"661c11fc", -- 14c8
		x"0032fdd7", -- 14cc
		x"08380004", -- 14d0
		x"feda6606", -- 14d4
		x"11fc0031", -- 14d8
		x"fdd741f8", -- 14dc
		x"fdd26000", -- 14e0
		x"429c0838", -- 14e4
		x"0004feda", -- 14e8
		x"67f011fc", -- 14ec
		x"0033fdd7", -- 14f0
		x"60e82878", -- 14f4
		x"fed4197c", -- 14f8
		x"000100a9", -- 14fc
		x"197c001f", -- 1500
		x"00a87022", -- 1504
		x"6100392a", -- 1508
		x"08ac0002", -- 150c
		x"005c422c", -- 1510
		x"005d08ac", -- 1514
		x"0001005c", -- 1518
		x"08ac0005", -- 151c
		x"005c2a4f", -- 1520
		x"4dfa005c", -- 1524
		x"45f90042", -- 1528
		x"800347f9", -- 152c
		x"00428001", -- 1530
		x"082c0006", -- 1534
		x"000b6630", -- 1538
		x"203c0007", -- 153c
		x"a1206100", -- 1540
		x"4fc4663a", -- 1544
		x"720041f9", -- 1548
		x"00428003", -- 154c
		x"12107600", -- 1550
		x"141076ff", -- 1554
		x"b4016626", -- 1558
		x"c23c00f0", -- 155c
		x"0c010070", -- 1560
		x"661c0c00", -- 1564
		x"008e661a", -- 1568
		x"4a390047", -- 156c
		x"800508b8", -- 1570
		x"0003fed2", -- 1574
		x"41fa45d3", -- 1578
		x"61003902", -- 157c
		x"600c2e4d", -- 1580
		x"600841fa", -- 1584
		x"45c56100", -- 1588
		x"38f843f8", -- 158c
		x"fee070fa", -- 1590
		x"2878fed4", -- 1594
		x"082c0006", -- 1598
		x"000b671c", -- 159c
		x"b2fcff3a", -- 15a0
		x"6712b2fc", -- 15a4
		x"ff52670c", -- 15a8
		x"b2fcff58", -- 15ac
		x"6706b2fc", -- 15b0
		x"ffd06604", -- 15b4
		x"5c89600a", -- 15b8
		x"32fc4eb9", -- 15bc
		x"22fc0000", -- 15c0
		x"4db8b089", -- 15c4
		x"66ce0838", -- 15c8
		x"0003fed2", -- 15cc
		x"66066100", -- 15d0
		x"54d66004", -- 15d4
		x"610053c2", -- 15d8
		x"61005d14", -- 15dc
		x"610052d4", -- 15e0
		x"60004202", -- 15e4
		x"31fc4ef9", -- 15e8
		x"ffb821fc", -- 15ec
		x"00004dbe", -- 15f0
		x"ffba027c", -- 15f4
		x"f8ff4e75", -- 15f8
		x"2878fed4", -- 15fc
		x"082c0004", -- 1600
-- disable RAM preload
--		x"000b665c", -- 1604
		x"000b605c", -- 1604
		x"700f6100", -- 1608
		x"382841fa", -- 160c
		x"42de6100", -- 1610
		x"41b86100", -- 1614
		x"f878082c", -- 1618
		x"0000000a", -- 161c
		x"672c4dfa", -- 1620
		x"0024203c", -- 1624
		x"eeee1111", -- 1628
		x"22002401", -- 162c
		x"26022803", -- 1630
		x"2a042c05", -- 1634
		x"2e0641f8", -- 1638
		x"c00090fc", -- 163c
		x"002048d0", -- 1640
		x"00ff60f6", -- 1644
		x"d0fc0020", -- 1648
		x"60124dfa", -- 164c
		x"000e41f8", -- 1650
		x"c0005988", -- 1654
		x"20884e71", -- 1658
		x"60f85888", -- 165c
		x"29480330", -- 1660
		x"6100f808", -- 1664
		x"41fa432e", -- 1668
		x"6100415e", -- 166c
		x"4e75702f", -- 1670
		x"610037be", -- 1674
		x"76ff78ff", -- 1678
		x"4dfa00d8", -- 167c
		x"2a4f0838", -- 1680
		x"0004fed2", -- 1684
		x"676245f9", -- 1688
		x"00520000", -- 168c
		x"43f90054", -- 1690
		x"00000839", -- 1694
		x"00040051", -- 1698
		x"fffe660a", -- 169c
		x"08390003", -- 16a0
		x"0051fffe", -- 16a4
		x"67420839", -- 16a8
		x"00030051", -- 16ac
		x"fffe6744", -- 16b0
		x"43f90056", -- 16b4
		x"00000839", -- 16b8
		x"00040051", -- 16bc
		x"fffe6634", -- 16c0
		x"264a2849", -- 16c4
		x"2e3c0f0f", -- 16c8
		x"0f0f6100", -- 16cc
		x"38364a40", -- 16d0
		x"6638244b", -- 16d4
		x"224c524a", -- 16d8
		x"52494dfa", -- 16dc
		x"00766100", -- 16e0
		x"38224a40", -- 16e4
		x"6624603c", -- 16e8
		x"45f90053", -- 16ec
		x"800043f9", -- 16f0
		x"00540000", -- 16f4
		x"08380001", -- 16f8
		x"fed2661c", -- 16fc
		x"524a5249", -- 1700
		x"7eff6100", -- 1704
		x"37fe4a40", -- 1708
		x"671a41fa", -- 170c
		x"44736100", -- 1710
		x"37706100", -- 1714
		x"39066038", -- 1718
		x"4a522a4a", -- 171c
		x"6100386c", -- 1720
		x"4a0066e6", -- 1724
		x"08380004", -- 1728
		x"fed26718", -- 172c
		x"41fa4442", -- 1730
		x"08390004", -- 1734
		x"0051fffe", -- 1738
		x"660e0839", -- 173c
		x"00030051", -- 1740
		x"fffe6604", -- 1744
		x"41fa4439", -- 1748
		x"61003732", -- 174c
		x"61003efe", -- 1750
		x"4e752e4d", -- 1754
		x"4e7550f8", -- 1758
		x"fed84e75", -- 175c
		x"4dfa0016", -- 1760
		x"1039005d", -- 1764
		x"00010c00", -- 1768
		x"002a6608", -- 176c
		x"41fa4474", -- 1770
		x"6100370a", -- 1774
		x"4e757028", -- 1778
		x"610036b6", -- 177c
		x"2878fed4", -- 1780
		x"422c033f", -- 1784
		x"4dfa007c", -- 1788
		x"4a790050", -- 178c
		x"00002878", -- 1790
		x"fed408ec", -- 1794
		x"0005000b", -- 1798
		x"323c2042", -- 179c
		x"197c0002", -- 17a0
		x"033f4dfa", -- 17a4
		x"00184a79", -- 17a8
		x"00508000", -- 17ac
		x"323c2041", -- 17b0
		x"197c0001", -- 17b4
		x"033f41fa", -- 17b8
		x"43d6601c", -- 17bc
		x"4dfafff8", -- 17c0
		x"4a390050", -- 17c4
		x"0004197c", -- 17c8
		x"0003033f", -- 17cc
		x"32390050", -- 17d0
		x"0012e059", -- 17d4
		x"41fa43c0", -- 17d8
		x"43f8fdd2", -- 17dc
		x"6100330a", -- 17e0
		x"12c1e049", -- 17e4
		x"12c14eb9", -- 17e8
		x"00014f9a", -- 17ec
		x"670a08ac", -- 17f0
		x"0005000b", -- 17f4
		x"610003f2", -- 17f8
		x"421141f8", -- 17fc
		x"fdd26100", -- 1800
		x"367c4e75", -- 1804
		x"08380004", -- 1808
		x"feda6758", -- 180c
		x"00790040", -- 1810
		x"005f400e", -- 1814
		x"3f38ffc4", -- 1818
		x"2f38ffc6", -- 181c
		x"31fc4ef9", -- 1820
		x"ffc421fc", -- 1824
		x"00001894", -- 1828
		x"ffc641f8", -- 182c
		x"fdd2f280", -- 1830
		x"0000f310", -- 1834
		x"10280001", -- 1838
		x"41fa4380", -- 183c
		x"b03c0018", -- 1840
		x"670e41fa", -- 1844
		x"438ab03c", -- 1848
		x"00386704", -- 184c
		x"41fa435d", -- 1850
		x"6100362a", -- 1854
		x"0279ffbe", -- 1858
		x"005f400e", -- 185c
		x"21dfffc6", -- 1860
		x"31dfffc4", -- 1864
		x"4dfa0028", -- 1868
		x"1039005c", -- 186c
		x"00010200", -- 1870
		x"007f41fa", -- 1874
		x"43270c00", -- 1878
		x"000a670e", -- 187c
		x"41fa4325", -- 1880
		x"0c00004a", -- 1884
		x"670441fa", -- 1888
		x"43236100", -- 188c
		x"35f04e75", -- 1890
		x"2f7c0000", -- 1894
		x"18580002", -- 1898
		x"4e732878", -- 189c
		x"fed44eb9", -- 18a0
		x"00007c5e", -- 18a4
		x"4eba672c", -- 18a8
		x"08ac0003", -- 18ac
		x"000a45f9", -- 18b0
		x"00600000", -- 18b4
		x"4241b27c", -- 18b8
		x"00206c00", -- 18bc
		x"02ce4dfa", -- 18c0
		x"02c22a4f", -- 18c4
		x"2001082c", -- 18c8
		x"0003000a", -- 18cc
		x"6604807c", -- 18d0
		x"00406100", -- 18d4
		x"355c747f", -- 18d8
		x"c42a0001", -- 18dc
		x"2878fed4", -- 18e0
		x"0c410007", -- 18e4
		x"66080838", -- 18e8
		x"0005fed2", -- 18ec
		x"67046100", -- 18f0
		x"67106100", -- 18f4
		x"f1c46100", -- 18f8
		x"02fe76ff", -- 18fc
		x"78ffb5ec", -- 1900
		x"00a26700", -- 1904
		x"01f60c2c", -- 1908
		x"000400a6", -- 190c
		x"6610264a", -- 1910
		x"d7fc0000", -- 1914
		x"4000b7ec", -- 1918
		x"00a26700", -- 191c
		x"02a8b43c", -- 1920
		x"00096626", -- 1924
		x"08380003", -- 1928
		x"fed26700", -- 192c
		x"01ceb5ec", -- 1930
		x"00b26700", -- 1934
		x"020c082c", -- 1938
		x"0005005c", -- 193c
		x"670001bc", -- 1940
		x"08ac0005", -- 1944
		x"005c6000", -- 1948
		x"01f848e7", -- 194c
		x"80c0302c", -- 1950
		x"032e41f8", -- 1954
		x"fdd24211", -- 1958
		x"61003e22", -- 195c
		x"3940032e", -- 1960
		x"4cdf0301", -- 1964
		x"b43c0034", -- 1968
		x"66160c2a", -- 196c
		x"00014001", -- 1970
		x"6600017e", -- 1974
		x"102a400d", -- 1978
		x"670001b8", -- 197c
		x"60000172", -- 1980
		x"b43c0015", -- 1984
		x"660c4eba", -- 1988
		x"2e4248e7", -- 198c
		x"64646000", -- 1990
		x"01581002", -- 1994
		x"0200001f", -- 1998
		x"0c000007", -- 199c
		x"66144219", -- 19a0
		x"41f8fdd2", -- 19a4
		x"4eba3dd6", -- 19a8
		x"4eb90001", -- 19ac
		x"67426000", -- 19b0
		x"0174b43c", -- 19b4
		x"00516618", -- 19b8
		x"082a0005", -- 19bc
		x"00056700", -- 19c0
		x"0130082a", -- 19c4
		x"00040005", -- 19c8
		x"66000126", -- 19cc
		x"60000164", -- 19d0
		x"b43c001c", -- 19d4
		x"660c48e7", -- 19d8
		x"64646100", -- 19dc
		x"305c6000", -- 19e0
		x"0108b43c", -- 19e4
		x"0001660c", -- 19e8
		x"48e76464", -- 19ec
		x"61002ee8", -- 19f0
		x"600000f6", -- 19f4
		x"b43c0008", -- 19f8
		x"660e4eb9", -- 19fc
		x"0001509e", -- 1a00
		x"67000130", -- 1a04
		x"600000ea", -- 1a08
		x"b43c0005", -- 1a0c
		x"662448e7", -- 1a10
		x"64646100", -- 1a14
		x"57f86000", -- 1a18
		x"00d02028", -- 1a1c
		x"436f6e73", -- 1a20
		x"6f6c6529", -- 1a24
		x"00202020", -- 1a28
		x"20747572", -- 1a2c
		x"6e206f6e", -- 1a30
		x"00002878", -- 1a34
		x"fed4b5ec", -- 1a38
		x"0048660c", -- 1a3c
		x"41faffdc", -- 1a40
		x"12d866fc", -- 1a44
		x"600000ec", -- 1a48
		x"1002c03c", -- 1a4c
		x"001f0c00", -- 1a50
		x"0019667e", -- 1a54
		x"082a0006", -- 1a58
		x"00016676", -- 1a5c
		x"421141f8", -- 1a60
		x"fdd26100", -- 1a64
		x"3d184dfa", -- 1a68
		x"001c4280", -- 1a6c
		x"010a0085", -- 1a70
		x"4a806710", -- 1a74
		x"4eb90000", -- 1a78
		x"7ce20838", -- 1a7c
		x"0005fdcc", -- 1a80
		x"660000a2", -- 1a84
		x"4dfa003e", -- 1a88
		x"43f8fdd2", -- 1a8c
		x"41faff97", -- 1a90
		x"12d866fc", -- 1a94
		x"53892a2c", -- 1a98
		x"004848e7", -- 1a9c
		x"e47c2a4f", -- 1aa0
		x"294a0048", -- 1aa4
		x"61003a66", -- 1aa8
		x"283c0000", -- 1aac
		x"4000204a", -- 1ab0
		x"61003424", -- 1ab4
		x"4cdf3e27", -- 1ab8
		x"29450048", -- 1abc
		x"4a436700", -- 1ac0
		x"0080600a", -- 1ac4
		x"2e4d4cdf", -- 1ac8
		x"3e272945", -- 1acc
		x"00482803", -- 1ad0
		x"601eb43c", -- 1ad4
		x"00026706", -- 1ad8
		x"b43c0042", -- 1adc
		x"661c5288", -- 1ae0
		x"48e76464", -- 1ae4
		x"61002ef2", -- 1ae8
		x"4cdf2626", -- 1aec
		x"4a00670a", -- 1af0
		x"610000f6", -- 1af4
		x"61006514", -- 1af8
		x"60382878", -- 1afc
		x"fed4082c", -- 1b00
		x"0003000a", -- 1b04
		x"672c4dfa", -- 1b08
		x"002a4280", -- 1b0c
		x"010a0085", -- 1b10
		x"4a80671e", -- 1b14
		x"421941f8", -- 1b18
		x"fdd26100", -- 1b1c
		x"3c604eb9", -- 1b20
		x"00007ce2", -- 1b24
		x"08380005", -- 1b28
		x"fdcc6714", -- 1b2c
		x"61003322", -- 1b30
		x"600e4219", -- 1b34
		x"41f8fdd2", -- 1b38
		x"61003c42", -- 1b3c
		x"610034dc", -- 1b40
		x"2878fed4", -- 1b44
		x"082c0003", -- 1b48
		x"000a6714", -- 1b4c
		x"42851a2a", -- 1b50
		x"0101e44d", -- 1b54
		x"5245d245", -- 1b58
		x"7416e5ad", -- 1b5c
		x"d5c56054", -- 1b60
		x"0c020051", -- 1b64
		x"671a7a1f", -- 1b68
		x"ca02ba3c", -- 1b6c
		x"001c6710", -- 1b70
		x"ba3c001d", -- 1b74
		x"670aba3c", -- 1b78
		x"001a6606", -- 1b7c
		x"615e615c", -- 1b80
		x"615a2e4d", -- 1b84
		x"61566000", -- 1b88
		x"fd2e2878", -- 1b8c
		x"fed4082c", -- 1b90
		x"0001000a", -- 1b94
		x"672c08ec", -- 1b98
		x"0003000a", -- 1b9c
		x"223c0000", -- 1ba0
		x"008445f9", -- 1ba4
		x"01000000", -- 1ba8
		x"60102e4d", -- 1bac
		x"d5fc0040", -- 1bb0
		x"00005241", -- 1bb4
		x"b27c0100", -- 1bb8
		x"6c084dfa", -- 1bbc
		x"ffee6000", -- 1bc0
		x"fd024e75", -- 1bc4
		x"0c2b000d", -- 1bc8
		x"4e476700", -- 1bcc
		x"ff240c2b", -- 1bd0
		x"000c4e47", -- 1bd4
		x"6700ff1a", -- 1bd8
		x"6000ff58", -- 1bdc
		x"5241d5fc", -- 1be0
		x"00010000", -- 1be4
		x"42824e75", -- 1be8
		x"61003266", -- 1bec
		x"41fa406a", -- 1bf0
		x"12d866fc", -- 1bf4
		x"4e7543f8", -- 1bf8
		x"fdd20c02", -- 1bfc
		x"00346600", -- 1c00
		x"00862878", -- 1c04
		x"fed46100", -- 1c08
		x"63ee674c", -- 1c0c
		x"707fc02a", -- 1c10
		x"0001b400", -- 1c14
		x"66420838", -- 1c18
		x"0001feda", -- 1c1c
		x"6628203c", -- 1c20
		x"004c4b40", -- 1c24
		x"2f004857", -- 1c28
		x"4eba35f0", -- 1c2c
		x"201f082a", -- 1c30
		x"00060003", -- 1c34
		x"66282f00", -- 1c38
		x"48574eba", -- 1c3c
		x"35fe6aec", -- 1c40
		x"588f7001", -- 1c44
		x"6006203c", -- 1c48
		x"000f4240", -- 1c4c
		x"082a0006", -- 1c50
		x"0003660a", -- 1c54
		x"53806ef4", -- 1c58
		x"41fa41f3", -- 1c5c
		x"603a0c2a", -- 1c60
		x"00014001", -- 1c64
		x"66f2102a", -- 1c68
		x"400d6706", -- 1c6c
		x"0c000006", -- 1c70
		x"66e641ea", -- 1c74
		x"400f32fc", -- 1c78
		x"48507005", -- 1c7c
		x"12d05448", -- 1c80
		x"53406ef8", -- 1c84
		x"602a41fa", -- 1c88
		x"401b1a18", -- 1c8c
		x"670aba02", -- 1c90
		x"67064a18", -- 1c94
		x"66fc60f2", -- 1c98
		x"12d866fc", -- 1c9c
		x"53894a05", -- 1ca0
		x"660e2002", -- 1ca4
		x"48e76000", -- 1ca8
		x"61002ddc", -- 1cac
		x"4cdf0006", -- 1cb0
		x"41fa3fa1", -- 1cb4
		x"12d866fc", -- 1cb8
		x"53894280", -- 1cbc
		x"100148e7", -- 1cc0
		x"60006100", -- 1cc4
		x"2dc24cdf", -- 1cc8
		x"0006204a", -- 1ccc
		x"4e757012", -- 1cd0
		x"6100315e", -- 1cd4
		x"2878fed4", -- 1cd8
		x"297c0002", -- 1cdc
		x"00000062", -- 1ce0
		x"197c005a", -- 1ce4
		x"006e244f", -- 1ce8
		x"4dfa00c8", -- 1cec
		x"206c0062", -- 1cf0
		x"b1fc0040", -- 1cf4
		x"00006400", -- 1cf8
		x"00c00c50", -- 1cfc
		x"f0ff660e", -- 1d00
		x"0c68f0ff", -- 1d04
		x"00026706", -- 1d08
		x"0c50f0ff", -- 1d0c
		x"670a06ac", -- 1d10
		x"00004000", -- 1d14
		x"006260d0", -- 1d18
		x"08280000", -- 1d1c
		x"00036706", -- 1d20
		x"19680002", -- 1d24
		x"006e1028", -- 1d28
		x"000c723f", -- 1d2c
		x"c0415240", -- 1d30
		x"c228000d", -- 1d34
		x"b0016660", -- 1d38
		x"08280000", -- 1d3c
		x"00036724", -- 1d40
		x"1028000e", -- 1d44
		x"08380000", -- 1d48
		x"fed26708", -- 1d4c
		x"08000006", -- 1d50
		x"67086010", -- 1d54
		x"08000003", -- 1d58
		x"660a2f08", -- 1d5c
		x"615c41fa", -- 1d60
		x"3eea603c", -- 1d64
		x"08280004", -- 1d68
		x"000366a2", -- 1d6c
		x"2f08283c", -- 1d70
		x"00004000", -- 1d74
		x"3028000e", -- 1d78
		x"0240f8f8", -- 1d7c
		x"0c404040", -- 1d80
		x"670a1028", -- 1d84
		x"00104880", -- 1d88
		x"e848c8c0", -- 1d8c
		x"61003118", -- 1d90
		x"205f4a40", -- 1d94
		x"6700ff78", -- 1d98
		x"2f08611e", -- 1d9c
		x"41fa3eba", -- 1da0
		x"12d866fc", -- 1da4
		x"41f8fdd2", -- 1da8
		x"610039d2", -- 1dac
		x"205f6000", -- 1db0
		x"ff5e2e4a", -- 1db4
		x"6000ff58", -- 1db8
		x"4e756100", -- 1dbc
		x"30942008", -- 1dc0
		x"43f8fdd2", -- 1dc4
		x"22fc524f", -- 1dc8
		x"4d2012ec", -- 1dcc
		x"006e41fa", -- 1dd0
		x"3e8312d8", -- 1dd4
		x"66fc5389", -- 1dd8
		x"60002cdc", -- 1ddc
		x"2878fed4", -- 1de0
		x"082c0004", -- 1de4
-- skip RAM test
		x"000b6600", -- 1de8
--		x"000b6000", -- 1de8
		x"00d4082c", -- 1dec
		x"0001000b", -- 1df0
		x"670000ca", -- 1df4
		x"70106100", -- 1df8
		x"303841fa", -- 1dfc
		x"3ade6100", -- 1e00
		x"39c808ac", -- 1e04
		x"0006000a", -- 1e08
		x"76ff78ff", -- 1e0c
		x"42b8fdd2", -- 1e10
		x"43f8ff22", -- 1e14
		x"32fc4ef9", -- 1e18
		x"22bc0000", -- 1e1c
		x"4c606100", -- 1e20
		x"f06c082c", -- 1e24
		x"0000000a", -- 1e28
		x"673243f8", -- 1e2c
		x"c0002a6c", -- 1e30
		x"0330487a", -- 1e34
		x"00124dfa", -- 1e38
		x"000a33fc", -- 1e3c
		x"0001005b", -- 1e40
		x"00006000", -- 1e44
		x"e8184dfa", -- 1e48
		x"00084279", -- 1e4c
		x"005b0000", -- 1e50
		x"2878fed4", -- 1e54
		x"266c0330", -- 1e58
		x"284d6052", -- 1e5c
		x"41ec0330", -- 1e60
		x"26504dfa", -- 1e64
		x"000a33fc", -- 1e68
		x"0001005b", -- 1e6c
		x"0000204b", -- 1e70
		x"284b5988", -- 1e74
		x"4dfa0022", -- 1e78
		x"600a4681", -- 1e7c
		x"2081b290", -- 1e80
		x"67f6600a", -- 1e84
		x"58882208", -- 1e88
		x"b2906612", -- 1e8c
		x"60ec2601", -- 1e90
		x"281049e8", -- 1e94
		x"000460e0", -- 1e98
		x"2848588c", -- 1e9c
		x"60dab0fc", -- 1ea0
		x"c00066ea", -- 1ea4
		x"4dfa0008", -- 1ea8
		x"4279005b", -- 1eac
		x"00006100", -- 1eb0
		x"efba2078", -- 1eb4
		x"fed408e8", -- 1eb8
		x"0006000a", -- 1ebc
		x"4e7541fa", -- 1ec0
		x"3ad46100", -- 1ec4
		x"39042078", -- 1ec8
		x"fed40828", -- 1ecc
		x"0004000b", -- 1ed0
		x"660000c8", -- 1ed4
		x"08280001", -- 1ed8
		x"000b6700", -- 1edc
		x"00542f0c", -- 1ee0
		x"b9cb673a", -- 1ee4
		x"61002f6a", -- 1ee8
		x"200c5980", -- 1eec
		x"21400328", -- 1ef0
		x"6100312c", -- 1ef4
		x"201f74ff", -- 1ef8
		x"42427601", -- 1efc
		x"4843b082", -- 1f00
		x"650c243c", -- 1f04
		x"fffff800", -- 1f08
		x"263c0000", -- 1f0c
		x"08002202", -- 1f10
		x"4681c280", -- 1f14
		x"6704c082", -- 1f18
		x"d0832f00", -- 1f1c
		x"601676ff", -- 1f20
		x"78ff6100", -- 1f24
		x"3182670c", -- 1f28
		x"70116100", -- 1f2c
		x"2f0460b4", -- 1f30
		x"2f280330", -- 1f34
		x"285f2078", -- 1f38
		x"fed4224c", -- 1f3c
		x"32280334", -- 1f40
		x"48c1eb89", -- 1f44
		x"d3c121c9", -- 1f48
		x"fdce40e7", -- 1f4c
		x"007c0700", -- 1f50
		x"2078fed4", -- 1f54
		x"224c323c", -- 1f58
		x"038812d8", -- 1f5c
		x"53416efa", -- 1f60
		x"21ccfed4", -- 1f64
		x"41ec00ca", -- 1f68
		x"294800b6", -- 1f6c
		x"08ec0004", -- 1f70
		x"000b46df", -- 1f74
		x"200cd0ac", -- 1f78
		x"002c4480", -- 1f7c
		x"43f8fdd2", -- 1f80
		x"22fc5241", -- 1f84
		x"4d206100", -- 1f88
		x"2afe41fa", -- 1f8c
		x"3c6a6100", -- 1f90
		x"2b5841f8", -- 1f94
		x"fdd26100", -- 1f98
		x"37e44e75", -- 1f9c
		x"ffffffff", -- 1fa0
		x"ffffffff", -- 1fa4
		x"ffffffff", -- 1fa8
		x"ffffffff", -- 1fac
		x"ffffffff", -- 1fb0
		x"ffffffff", -- 1fb4
		x"ffffffff", -- 1fb8
		x"ffffffff", -- 1fbc
		x"ffffffff", -- 1fc0
		x"ffffffff", -- 1fc4
		x"ffffffff", -- 1fc8
		x"ffffffff", -- 1fcc
		x"ffffffff", -- 1fd0
		x"ffffffff", -- 1fd4
		x"ffffffff", -- 1fd8
		x"ffffffff", -- 1fdc
		x"ffffffff", -- 1fe0
		x"ffffffff", -- 1fe4
		x"ffffffff", -- 1fe8
		x"ffffffff", -- 1fec
		x"ffffffff", -- 1ff0
		x"ffffffff", -- 1ff4
		x"ffffffff", -- 1ff8
		x"ffffffff", -- 1ffc
		x"00486858", -- 2000
		x"48001212", -- 2004
		x"121e0000", -- 2008
		x"00000000", -- 200c
		x"00384030", -- 2010
		x"08700012", -- 2014
		x"1e120000", -- 2018
		x"00000000", -- 201c
		x"00384030", -- 2020
		x"0870000a", -- 2024
		x"040a0000", -- 2028
		x"00000000", -- 202c
		x"00704060", -- 2030
		x"4070000a", -- 2034
		x"040a0000", -- 2038
		x"00000000", -- 203c
		x"00704060", -- 2040
		x"40700e04", -- 2044
		x"04040000", -- 2048
		x"00000000", -- 204c
		x"00704060", -- 2050
		x"40700c12", -- 2054
		x"160e0000", -- 2058
		x"00000000", -- 205c
		x"00304878", -- 2060
		x"48481014", -- 2064
		x"18140000", -- 2068
		x"00000000", -- 206c
		x"00081c22", -- 2070
		x"2222227f", -- 2074
		x"08080000", -- 2078
		x"00000000", -- 207c
		x"00704870", -- 2080
		x"48730402", -- 2084
		x"01060000", -- 2088
		x"00000000", -- 208c
		x"00484878", -- 2090
		x"48480702", -- 2094
		x"02020000", -- 2098
		x"00000000", -- 209c
		x"00404040", -- 20a0
		x"40770406", -- 20a4
		x"04040000", -- 20a8
		x"00000000", -- 20ac
		x"00444428", -- 20b0
		x"10000e04", -- 20b4
		x"04040000", -- 20b8
		x"00000000", -- 20bc
		x"00784070", -- 20c0
		x"404f080e", -- 20c4
		x"08080000", -- 20c8
		x"00000000", -- 20cc
		x"00384040", -- 20d0
		x"380e090e", -- 20d4
		x"0a090000", -- 20d8
		x"00000000", -- 20dc
		x"00384030", -- 20e0
		x"08760909", -- 20e4
		x"09060000", -- 20e8
		x"00000000", -- 20ec
		x"00384030", -- 20f0
		x"08770202", -- 20f4
		x"02070000", -- 20f8
		x"00000000", -- 20fc
		x"00704848", -- 2100
		x"48700404", -- 2104
		x"04070000", -- 2108
		x"00000000", -- 210c
		x"00704848", -- 2110
		x"48720602", -- 2114
		x"02070000", -- 2118
		x"00000000", -- 211c
		x"00704848", -- 2120
		x"48760102", -- 2124
		x"04070000", -- 2128
		x"00000000", -- 212c
		x"00704848", -- 2130
		x"48770103", -- 2134
		x"01070000", -- 2138
		x"00000000", -- 213c
		x"00704848", -- 2140
		x"4872060f", -- 2144
		x"02020000", -- 2148
		x"00000000", -- 214c
		x"00486858", -- 2150
		x"48040506", -- 2154
		x"06050000", -- 2158
		x"00000000", -- 215c
		x"00384030", -- 2160
		x"08700502", -- 2164
		x"02020000", -- 2168
		x"00000000", -- 216c
		x"00704060", -- 2170
		x"40760506", -- 2174
		x"05060000", -- 2178
		x"00000000", -- 217c
		x"00384040", -- 2180
		x"3800090d", -- 2184
		x"0b090000", -- 2188
		x"00000000", -- 218c
		x"00784060", -- 2190
		x"4078111b", -- 2194
		x"15110000", -- 2198
		x"00000000", -- 219c
		x"00384030", -- 21a0
		x"08760506", -- 21a4
		x"05060000", -- 21a8
		x"00000000", -- 21ac
		x"00784070", -- 21b0
		x"40780304", -- 21b4
		x"04030000", -- 21b8
		x"00000000", -- 21bc
		x"00784070", -- 21c0
		x"40470806", -- 21c4
		x"010e0000", -- 21c8
		x"00000000", -- 21cc
		x"00384058", -- 21d0
		x"483f0806", -- 21d4
		x"010e0000", -- 21d8
		x"00000000", -- 21dc
		x"00704870", -- 21e0
		x"50570806", -- 21e4
		x"010e0000", -- 21e8
		x"00000000", -- 21ec
		x"00484848", -- 21f0
		x"78070806", -- 21f4
		x"010e0000", -- 21f8
		x"00000000", -- 21fc
		x"00000000", -- 2200
		x"00000000", -- 2204
		x"00000000", -- 2208
		x"00000000", -- 220c
		x"00101010", -- 2210
		x"10100010", -- 2214
		x"00000000", -- 2218
		x"00000000", -- 221c
		x"00282828", -- 2220
		x"00000000", -- 2224
		x"00000000", -- 2228
		x"00000000", -- 222c
		x"0028287c", -- 2230
		x"287c2828", -- 2234
		x"00000000", -- 2238
		x"00000000", -- 223c
		x"00103c50", -- 2240
		x"38147810", -- 2244
		x"00000000", -- 2248
		x"00000000", -- 224c
		x"00606408", -- 2250
		x"10204c0c", -- 2254
		x"00000000", -- 2258
		x"00000000", -- 225c
		x"00205050", -- 2260
		x"20544834", -- 2264
		x"00000000", -- 2268
		x"00000000", -- 226c
		x"00081020", -- 2270
		x"00000000", -- 2274
		x"00000000", -- 2278
		x"00000000", -- 227c
		x"00081010", -- 2280
		x"10101008", -- 2284
		x"00000000", -- 2288
		x"00000000", -- 228c
		x"00100808", -- 2290
		x"08080810", -- 2294
		x"00000000", -- 2298
		x"00000000", -- 229c
		x"00002810", -- 22a0
		x"7c102800", -- 22a4
		x"00000000", -- 22a8
		x"00000000", -- 22ac
		x"00001010", -- 22b0
		x"7c101000", -- 22b4
		x"00000000", -- 22b8
		x"00000000", -- 22bc
		x"00000000", -- 22c0
		x"00001818", -- 22c4
		x"08100000", -- 22c8
		x"00000000", -- 22cc
		x"00000000", -- 22d0
		x"7c000000", -- 22d4
		x"00000000", -- 22d8
		x"00000000", -- 22dc
		x"00000000", -- 22e0
		x"00001818", -- 22e4
		x"00000000", -- 22e8
		x"00000000", -- 22ec
		x"00000408", -- 22f0
		x"10204000", -- 22f4
		x"00000000", -- 22f8
		x"00000000", -- 22fc
		x"0038444c", -- 2300
		x"54644438", -- 2304
		x"00000000", -- 2308
		x"00000000", -- 230c
		x"00103010", -- 2310
		x"10101038", -- 2314
		x"00000000", -- 2318
		x"00000000", -- 231c
		x"00384404", -- 2320
		x"0830407c", -- 2324
		x"00000000", -- 2328
		x"00000000", -- 232c
		x"00384404", -- 2330
		x"18044438", -- 2334
		x"00000000", -- 2338
		x"00000000", -- 233c
		x"00081828", -- 2340
		x"487c0808", -- 2344
		x"00000000", -- 2348
		x"00000000", -- 234c
		x"007c4078", -- 2350
		x"04044438", -- 2354
		x"00000000", -- 2358
		x"00000000", -- 235c
		x"001c2040", -- 2360
		x"78444438", -- 2364
		x"00000000", -- 2368
		x"00000000", -- 236c
		x"007c0408", -- 2370
		x"10202020", -- 2374
		x"00000000", -- 2378
		x"00000000", -- 237c
		x"00384444", -- 2380
		x"38444438", -- 2384
		x"00000000", -- 2388
		x"00000000", -- 238c
		x"00384444", -- 2390
		x"3c040830", -- 2394
		x"00000000", -- 2398
		x"00000000", -- 239c
		x"00001818", -- 23a0
		x"00001818", -- 23a4
		x"00000000", -- 23a8
		x"00000000", -- 23ac
		x"00001818", -- 23b0
		x"00001818", -- 23b4
		x"08100000", -- 23b8
		x"00000000", -- 23bc
		x"00081020", -- 23c0
		x"40201008", -- 23c4
		x"00000000", -- 23c8
		x"00000000", -- 23cc
		x"0000007c", -- 23d0
		x"007c0000", -- 23d4
		x"00000000", -- 23d8
		x"00000000", -- 23dc
		x"00201008", -- 23e0
		x"04081020", -- 23e4
		x"00000000", -- 23e8
		x"00000000", -- 23ec
		x"00384404", -- 23f0
		x"08100010", -- 23f4
		x"00000000", -- 23f8
		x"00000000", -- 23fc
		x"0038445c", -- 2400
		x"545c4038", -- 2404
		x"00000000", -- 2408
		x"00000000", -- 240c
		x"00384444", -- 2410
		x"7c444444", -- 2414
		x"00000000", -- 2418
		x"00000000", -- 241c
		x"00782424", -- 2420
		x"38242478", -- 2424
		x"00000000", -- 2428
		x"00000000", -- 242c
		x"00384440", -- 2430
		x"40404438", -- 2434
		x"00000000", -- 2438
		x"00000000", -- 243c
		x"00782424", -- 2440
		x"24242478", -- 2444
		x"00000000", -- 2448
		x"00000000", -- 244c
		x"007c4040", -- 2450
		x"7840407c", -- 2454
		x"00000000", -- 2458
		x"00000000", -- 245c
		x"007c4040", -- 2460
		x"78404040", -- 2464
		x"00000000", -- 2468
		x"00000000", -- 246c
		x"00384440", -- 2470
		x"404c4438", -- 2474
		x"00000000", -- 2478
		x"00000000", -- 247c
		x"00444444", -- 2480
		x"7c444444", -- 2484
		x"00000000", -- 2488
		x"00000000", -- 248c
		x"00381010", -- 2490
		x"10101038", -- 2494
		x"00000000", -- 2498
		x"00000000", -- 249c
		x"001c0808", -- 24a0
		x"08084830", -- 24a4
		x"00000000", -- 24a8
		x"00000000", -- 24ac
		x"00444850", -- 24b0
		x"60504844", -- 24b4
		x"00000000", -- 24b8
		x"00000000", -- 24bc
		x"00404040", -- 24c0
		x"4040407c", -- 24c4
		x"00000000", -- 24c8
		x"00000000", -- 24cc
		x"00446c54", -- 24d0
		x"54444444", -- 24d4
		x"00000000", -- 24d8
		x"00000000", -- 24dc
		x"00444464", -- 24e0
		x"544c4444", -- 24e4
		x"00000000", -- 24e8
		x"00000000", -- 24ec
		x"00384444", -- 24f0
		x"44444438", -- 24f4
		x"00000000", -- 24f8
		x"00000000", -- 24fc
		x"00784444", -- 2500
		x"78404040", -- 2504
		x"00000000", -- 2508
		x"00000000", -- 250c
		x"00384444", -- 2510
		x"44544834", -- 2514
		x"00000000", -- 2518
		x"00000000", -- 251c
		x"00784444", -- 2520
		x"78504844", -- 2524
		x"00000000", -- 2528
		x"00000000", -- 252c
		x"00384440", -- 2530
		x"38044438", -- 2534
		x"00000000", -- 2538
		x"00000000", -- 253c
		x"007c1010", -- 2540
		x"10101010", -- 2544
		x"00000000", -- 2548
		x"00000000", -- 254c
		x"00444444", -- 2550
		x"44444438", -- 2554
		x"00000000", -- 2558
		x"00000000", -- 255c
		x"00444444", -- 2560
		x"28281010", -- 2564
		x"00000000", -- 2568
		x"00000000", -- 256c
		x"00444444", -- 2570
		x"54546c44", -- 2574
		x"00000000", -- 2578
		x"00000000", -- 257c
		x"00444428", -- 2580
		x"10284444", -- 2584
		x"00000000", -- 2588
		x"00000000", -- 258c
		x"00444428", -- 2590
		x"10101010", -- 2594
		x"00000000", -- 2598
		x"00000000", -- 259c
		x"007c0408", -- 25a0
		x"1020407c", -- 25a4
		x"00000000", -- 25a8
		x"00000000", -- 25ac
		x"00382020", -- 25b0
		x"20202038", -- 25b4
		x"00000000", -- 25b8
		x"00000000", -- 25bc
		x"00004020", -- 25c0
		x"10080400", -- 25c4
		x"00000000", -- 25c8
		x"00000000", -- 25cc
		x"00380808", -- 25d0
		x"08080838", -- 25d4
		x"00000000", -- 25d8
		x"00000000", -- 25dc
		x"00102844", -- 25e0
		x"00000000", -- 25e4
		x"00000000", -- 25e8
		x"00000000", -- 25ec
		x"00000000", -- 25f0
		x"00000000", -- 25f4
		x"00ff0000", -- 25f8
		x"00000000", -- 25fc
		x"00201008", -- 2600
		x"00000000", -- 2604
		x"00000000", -- 2608
		x"00000000", -- 260c
		x"00000038", -- 2610
		x"043c443e", -- 2614
		x"00000000", -- 2618
		x"00000000", -- 261c
		x"00404078", -- 2620
		x"44444478", -- 2624
		x"00000000", -- 2628
		x"00000000", -- 262c
		x"00000038", -- 2630
		x"40404038", -- 2634
		x"00000000", -- 2638
		x"00000000", -- 263c
		x"0004043c", -- 2640
		x"4444443c", -- 2644
		x"00000000", -- 2648
		x"00000000", -- 264c
		x"00000038", -- 2650
		x"44784038", -- 2654
		x"00000000", -- 2658
		x"00000000", -- 265c
		x"00182420", -- 2660
		x"70202020", -- 2664
		x"00000000", -- 2668
		x"00000000", -- 266c
		x"0000003c", -- 2670
		x"4444443c", -- 2674
		x"04443800", -- 2678
		x"00000000", -- 267c
		x"00404058", -- 2680
		x"64444444", -- 2684
		x"00000000", -- 2688
		x"00000000", -- 268c
		x"00100030", -- 2690
		x"10101010", -- 2694
		x"00000000", -- 2698
		x"00000000", -- 269c
		x"00080018", -- 26a0
		x"08080808", -- 26a4
		x"48300000", -- 26a8
		x"00000000", -- 26ac
		x"00202024", -- 26b0
		x"28302824", -- 26b4
		x"00000000", -- 26b8
		x"00000000", -- 26bc
		x"00180808", -- 26c0
		x"08080808", -- 26c4
		x"00000000", -- 26c8
		x"00000000", -- 26cc
		x"00000068", -- 26d0
		x"54545454", -- 26d4
		x"00000000", -- 26d8
		x"00000000", -- 26dc
		x"00000058", -- 26e0
		x"64444444", -- 26e4
		x"00000000", -- 26e8
		x"00000000", -- 26ec
		x"00000038", -- 26f0
		x"44444438", -- 26f4
		x"00000000", -- 26f8
		x"00000000", -- 26fc
		x"00000058", -- 2700
		x"64446458", -- 2704
		x"40404000", -- 2708
		x"00000000", -- 270c
		x"00000034", -- 2710
		x"4c444c34", -- 2714
		x"04040400", -- 2718
		x"00000000", -- 271c
		x"00000058", -- 2720
		x"64404040", -- 2724
		x"00000000", -- 2728
		x"00000000", -- 272c
		x"00000038", -- 2730
		x"40380478", -- 2734
		x"00000000", -- 2738
		x"00000000", -- 273c
		x"00202070", -- 2740
		x"20202810", -- 2744
		x"00000000", -- 2748
		x"00000000", -- 274c
		x"00000044", -- 2750
		x"44444c34", -- 2754
		x"00000000", -- 2758
		x"00000000", -- 275c
		x"00000044", -- 2760
		x"44442810", -- 2764
		x"00000000", -- 2768
		x"00000000", -- 276c
		x"00000044", -- 2770
		x"54545428", -- 2774
		x"00000000", -- 2778
		x"00000000", -- 277c
		x"00000044", -- 2780
		x"28102844", -- 2784
		x"00000000", -- 2788
		x"00000000", -- 278c
		x"00000044", -- 2790
		x"44442818", -- 2794
		x"10204000", -- 2798
		x"00000000", -- 279c
		x"0000007c", -- 27a0
		x"0810207c", -- 27a4
		x"00000000", -- 27a8
		x"00000000", -- 27ac
		x"08101010", -- 27b0
		x"20101010", -- 27b4
		x"08000000", -- 27b8
		x"00000000", -- 27bc
		x"10101010", -- 27c0
		x"10101010", -- 27c4
		x"10101010", -- 27c8
		x"00000000", -- 27cc
		x"20101010", -- 27d0
		x"08101010", -- 27d4
		x"20000000", -- 27d8
		x"00000000", -- 27dc
		x"00000000", -- 27e0
		x"20540800", -- 27e4
		x"00000000", -- 27e8
		x"00000000", -- 27ec
		x"00285428", -- 27f0
		x"54285428", -- 27f4
		x"00000000", -- 27f8
		x"00000000", -- 27fc
		x"0044287c", -- 2800
		x"107c1010", -- 2804
		x"00000000", -- 2808
		x"00000000", -- 280c
		x"00000000", -- 2810
		x"30484830", -- 2814
		x"00000000", -- 2818
		x"00000000", -- 281c
		x"001c1010", -- 2820
		x"10000000", -- 2824
		x"00000000", -- 2828
		x"00000000", -- 282c
		x"00000000", -- 2830
		x"10101070", -- 2834
		x"00000000", -- 2838
		x"00000000", -- 283c
		x"00000000", -- 2840
		x"00402010", -- 2844
		x"00000000", -- 2848
		x"00000000", -- 284c
		x"00000000", -- 2850
		x"30300000", -- 2854
		x"00000000", -- 2858
		x"00000000", -- 285c
		x"00007c04", -- 2860
		x"7c040810", -- 2864
		x"00000000", -- 2868
		x"00000000", -- 286c
		x"0000007c", -- 2870
		x"04181020", -- 2874
		x"00000000", -- 2878
		x"00000000", -- 287c
		x"00000008", -- 2880
		x"10305010", -- 2884
		x"00000000", -- 2888
		x"00000000", -- 288c
		x"00000010", -- 2890
		x"7c440418", -- 2894
		x"00000000", -- 2898
		x"00000000", -- 289c
		x"00000000", -- 28a0
		x"7c10107c", -- 28a4
		x"00000000", -- 28a8
		x"00000000", -- 28ac
		x"00000008", -- 28b0
		x"7c182848", -- 28b4
		x"00000000", -- 28b8
		x"00000000", -- 28bc
		x"00000020", -- 28c0
		x"7c242820", -- 28c4
		x"00000000", -- 28c8
		x"00000000", -- 28cc
		x"00000000", -- 28d0
		x"3808087c", -- 28d4
		x"00000000", -- 28d8
		x"00000000", -- 28dc
		x"00000078", -- 28e0
		x"08780878", -- 28e4
		x"00000000", -- 28e8
		x"00000000", -- 28ec
		x"00000000", -- 28f0
		x"54540418", -- 28f4
		x"00000000", -- 28f8
		x"00000000", -- 28fc
		x"00000000", -- 2900
		x"7c000000", -- 2904
		x"00000000", -- 2908
		x"00000000", -- 290c
		x"007c0414", -- 2910
		x"18101020", -- 2914
		x"00000000", -- 2918
		x"00000000", -- 291c
		x"00040810", -- 2920
		x"30501010", -- 2924
		x"00000000", -- 2928
		x"00000000", -- 292c
		x"00107c44", -- 2930
		x"44040810", -- 2934
		x"00000000", -- 2938
		x"00000000", -- 293c
		x"00007c10", -- 2940
		x"1010107c", -- 2944
		x"00000000", -- 2948
		x"00000000", -- 294c
		x"00087c08", -- 2950
		x"18284808", -- 2954
		x"00000000", -- 2958
		x"00000000", -- 295c
		x"00207c24", -- 2960
		x"24242448", -- 2964
		x"00000000", -- 2968
		x"00000000", -- 296c
		x"00107c10", -- 2970
		x"7c101010", -- 2974
		x"00000000", -- 2978
		x"00000000", -- 297c
		x"00003c24", -- 2980
		x"44040830", -- 2984
		x"00000000", -- 2988
		x"00000000", -- 298c
		x"00203c48", -- 2990
		x"08080810", -- 2994
		x"00000000", -- 2998
		x"00000000", -- 299c
		x"00007c04", -- 29a0
		x"0404047c", -- 29a4
		x"00000000", -- 29a8
		x"00000000", -- 29ac
		x"00287c28", -- 29b0
		x"28081020", -- 29b4
		x"00000000", -- 29b8
		x"00000000", -- 29bc
		x"00006004", -- 29c0
		x"64040870", -- 29c4
		x"00000000", -- 29c8
		x"00000000", -- 29cc
		x"00007c04", -- 29d0
		x"08102844", -- 29d4
		x"00000000", -- 29d8
		x"00000000", -- 29dc
		x"00207c24", -- 29e0
		x"2820201c", -- 29e4
		x"00000000", -- 29e8
		x"00000000", -- 29ec
		x"00004444", -- 29f0
		x"24040830", -- 29f4
		x"00000000", -- 29f8
		x"00000000", -- 29fc
		x"00003c24", -- 2a00
		x"540c0830", -- 2a04
		x"00000000", -- 2a08
		x"00000000", -- 2a0c
		x"00087010", -- 2a10
		x"7c101020", -- 2a14
		x"00000000", -- 2a18
		x"00000000", -- 2a1c
		x"00005454", -- 2a20
		x"54040810", -- 2a24
		x"00000000", -- 2a28
		x"00000000", -- 2a2c
		x"0038007c", -- 2a30
		x"10101020", -- 2a34
		x"00000000", -- 2a38
		x"00000000", -- 2a3c
		x"00202020", -- 2a40
		x"30282020", -- 2a44
		x"00000000", -- 2a48
		x"00000000", -- 2a4c
		x"0010107c", -- 2a50
		x"10101020", -- 2a54
		x"00000000", -- 2a58
		x"00000000", -- 2a5c
		x"00003800", -- 2a60
		x"0000007c", -- 2a64
		x"00000000", -- 2a68
		x"00000000", -- 2a6c
		x"00007c04", -- 2a70
		x"28102840", -- 2a74
		x"00000000", -- 2a78
		x"00000000", -- 2a7c
		x"08100000", -- 2a80
		x"00000000", -- 2a84
		x"00000000", -- 2a88
		x"00000000", -- 2a8c
		x"20100000", -- 2a90
		x"00000000", -- 2a94
		x"00000000", -- 2a98
		x"00000000", -- 2a9c
		x"10280000", -- 2aa0
		x"00000000", -- 2aa4
		x"00000000", -- 2aa8
		x"00000000", -- 2aac
		x"00280000", -- 2ab0
		x"00000000", -- 2ab4
		x"00000000", -- 2ab8
		x"00000000", -- 2abc
		x"20540800", -- 2ac0
		x"00000000", -- 2ac4
		x"00000000", -- 2ac8
		x"00000000", -- 2acc
		x"00107c08", -- 2ad0
		x"10385410", -- 2ad4
		x"00000000", -- 2ad8
		x"00000000", -- 2adc
		x"00080808", -- 2ae0
		x"08081020", -- 2ae4
		x"00000000", -- 2ae8
		x"00000000", -- 2aec
		x"1c222070", -- 2af0
		x"20702022", -- 2af4
		x"7c000000", -- 2af8
		x"00000000", -- 2afc
		x"ff000000", -- 2b00
		x"00000000", -- 2b04
		x"00000000", -- 2b08
		x"00000000", -- 2b0c
		x"00001008", -- 2b10
		x"44444444", -- 2b14
		x"00000000", -- 2b18
		x"00000000", -- 2b1c
		x"0040407c", -- 2b20
		x"4040403c", -- 2b24
		x"00000000", -- 2b28
		x"00000000", -- 2b2c
		x"30484830", -- 2b30
		x"00000000", -- 2b34
		x"00000000", -- 2b38
		x"00000000", -- 2b3c
		x"00007c04", -- 2b40
		x"04040830", -- 2b44
		x"00000000", -- 2b48
		x"00000000", -- 2b4c
		x"00000038", -- 2b50
		x"40404438", -- 2b54
		x"10083000", -- 2b58
		x"00000000", -- 2b5c
		x"20540844", -- 2b60
		x"64544c44", -- 2b64
		x"00000000", -- 2b68
		x"00000000", -- 2b6c
		x"20540800", -- 2b70
		x"58644444", -- 2b74
		x"00000000", -- 2b78
		x"00000000", -- 2b7c
		x"00100010", -- 2b80
		x"10101010", -- 2b84
		x"00000000", -- 2b88
		x"00000000", -- 2b8c
		x"00100010", -- 2b90
		x"20404438", -- 2b94
		x"00000000", -- 2b98
		x"00000000", -- 2b9c
		x"0000423c", -- 2ba0
		x"24243c42", -- 2ba4
		x"00000000", -- 2ba8
		x"00000000", -- 2bac
		x"1c222020", -- 2bb0
		x"7020227c", -- 2bb4
		x"00000000", -- 2bb8
		x"00000000", -- 2bbc
		x"00002050", -- 2bc0
		x"08040400", -- 2bc4
		x"00000000", -- 2bc8
		x"00000000", -- 2bcc
		x"18242010", -- 2bd0
		x"38241c08", -- 2bd4
		x"04241800", -- 2bd8
		x"00000000", -- 2bdc
		x"00107c10", -- 2be0
		x"54545410", -- 2be4
		x"00000000", -- 2be8
		x"00000000", -- 2bec
		x"00007c04", -- 2bf0
		x"04281008", -- 2bf4
		x"00000000", -- 2bf8
		x"00000000", -- 2bfc
		x"10280038", -- 2c00
		x"043c443e", -- 2c04
		x"00000000", -- 2c08
		x"00000000", -- 2c0c
		x"10280038", -- 2c10
		x"44784038", -- 2c14
		x"00000000", -- 2c18
		x"00000000", -- 2c1c
		x"10280038", -- 2c20
		x"44444438", -- 2c24
		x"00000000", -- 2c28
		x"00000000", -- 2c2c
		x"10280044", -- 2c30
		x"44444c34", -- 2c34
		x"00000000", -- 2c38
		x"00000000", -- 2c3c
		x"08100038", -- 2c40
		x"043c443e", -- 2c44
		x"00000000", -- 2c48
		x"00000000", -- 2c4c
		x"08100038", -- 2c50
		x"44784038", -- 2c54
		x"00000000", -- 2c58
		x"00000000", -- 2c5c
		x"08100038", -- 2c60
		x"44444438", -- 2c64
		x"00000000", -- 2c68
		x"00000000", -- 2c6c
		x"08100044", -- 2c70
		x"44444c34", -- 2c74
		x"00000000", -- 2c78
		x"00000000", -- 2c7c
		x"20100038", -- 2c80
		x"043c443e", -- 2c84
		x"00000000", -- 2c88
		x"00000000", -- 2c8c
		x"20100038", -- 2c90
		x"44784038", -- 2c94
		x"00000000", -- 2c98
		x"00000000", -- 2c9c
		x"20100038", -- 2ca0
		x"44444438", -- 2ca4
		x"00000000", -- 2ca8
		x"00000000", -- 2cac
		x"20100044", -- 2cb0
		x"44444c34", -- 2cb4
		x"00000000", -- 2cb8
		x"00000000", -- 2cbc
		x"00280038", -- 2cc0
		x"043c443e", -- 2cc4
		x"00000000", -- 2cc8
		x"00000000", -- 2ccc
		x"00280038", -- 2cd0
		x"44784038", -- 2cd4
		x"00000000", -- 2cd8
		x"00000000", -- 2cdc
		x"00280038", -- 2ce0
		x"44444438", -- 2ce4
		x"00000000", -- 2ce8
		x"00000000", -- 2cec
		x"00280044", -- 2cf0
		x"44444c34", -- 2cf4
		x"00000000", -- 2cf8
		x"00000000", -- 2cfc
		x"10003844", -- 2d00
		x"447c4444", -- 2d04
		x"00000000", -- 2d08
		x"00000000", -- 2d0c
		x"10280010", -- 2d10
		x"10101010", -- 2d14
		x"00000000", -- 2d18
		x"00000000", -- 2d1c
		x"003c4c4c", -- 2d20
		x"54646478", -- 2d24
		x"00000000", -- 2d28
		x"00000000", -- 2d2c
		x"003e5090", -- 2d30
		x"fc90909e", -- 2d34
		x"00000000", -- 2d38
		x"00000000", -- 2d3c
		x"00100038", -- 2d40
		x"043c443e", -- 2d44
		x"00000000", -- 2d48
		x"00000000", -- 2d4c
		x"08100010", -- 2d50
		x"10101010", -- 2d54
		x"00000000", -- 2d58
		x"00000000", -- 2d5c
		x"0000003c", -- 2d60
		x"4c546478", -- 2d64
		x"00000000", -- 2d68
		x"00000000", -- 2d6c
		x"000000ec", -- 2d70
		x"127c906e", -- 2d74
		x"00000000", -- 2d78
		x"00000000", -- 2d7c
		x"28003844", -- 2d80
		x"447c4444", -- 2d84
		x"00000000", -- 2d88
		x"00000000", -- 2d8c
		x"20100010", -- 2d90
		x"10101010", -- 2d94
		x"00000000", -- 2d98
		x"00000000", -- 2d9c
		x"28003844", -- 2da0
		x"44444438", -- 2da4
		x"00000000", -- 2da8
		x"00000000", -- 2dac
		x"28004444", -- 2db0
		x"44444438", -- 2db4
		x"00000000", -- 2db8
		x"00000000", -- 2dbc
		x"08107c40", -- 2dc0
		x"7040407c", -- 2dc4
		x"00000000", -- 2dc8
		x"00000000", -- 2dcc
		x"00280010", -- 2dd0
		x"10101010", -- 2dd4
		x"00000000", -- 2dd8
		x"00000000", -- 2ddc
		x"00384444", -- 2de0
		x"58444458", -- 2de4
		x"40000000", -- 2de8
		x"00000000", -- 2dec
		x"00404060", -- 2df0
		x"50500c0a", -- 2df4
		x"0c080800", -- 2df8
		x"00000000", -- 2dfc
		x"00003800", -- 2e00
		x"38003804", -- 2e04
		x"00000000", -- 2e08
		x"00000000", -- 2e0c
		x"00001020", -- 2e10
		x"40447c04", -- 2e14
		x"00000000", -- 2e18
		x"00000000", -- 2e1c
		x"00000404", -- 2e20
		x"28102840", -- 2e24
		x"00000000", -- 2e28
		x"00000000", -- 2e2c
		x"00007c20", -- 2e30
		x"7c20201c", -- 2e34
		x"00000000", -- 2e38
		x"00000000", -- 2e3c
		x"0020207c", -- 2e40
		x"24282020", -- 2e44
		x"00000000", -- 2e48
		x"00000000", -- 2e4c
		x"00003808", -- 2e50
		x"0808087c", -- 2e54
		x"00000000", -- 2e58
		x"00000000", -- 2e5c
		x"00007c04", -- 2e60
		x"7c04047c", -- 2e64
		x"00000000", -- 2e68
		x"00000000", -- 2e6c
		x"0038007c", -- 2e70
		x"04040810", -- 2e74
		x"00000000", -- 2e78
		x"00000000", -- 2e7c
		x"00484848", -- 2e80
		x"48081020", -- 2e84
		x"00000000", -- 2e88
		x"00000000", -- 2e8c
		x"00001050", -- 2e90
		x"50545458", -- 2e94
		x"00000000", -- 2e98
		x"00000000", -- 2e9c
		x"00004040", -- 2ea0
		x"44485060", -- 2ea4
		x"00000000", -- 2ea8
		x"00000000", -- 2eac
		x"00007c44", -- 2eb0
		x"4444447c", -- 2eb4
		x"00000000", -- 2eb8
		x"00000000", -- 2ebc
		x"00007c44", -- 2ec0
		x"44040810", -- 2ec4
		x"00000000", -- 2ec8
		x"00000000", -- 2ecc
		x"00006000", -- 2ed0
		x"04040870", -- 2ed4
		x"00000000", -- 2ed8
		x"00000000", -- 2edc
		x"00104820", -- 2ee0
		x"00000000", -- 2ee4
		x"00000000", -- 2ee8
		x"00000000", -- 2eec
		x"00001008", -- 2ef0
		x"7c081000", -- 2ef4
		x"00000000", -- 2ef8
		x"00000000", -- 2efc
		x"00003c20", -- 2f00
		x"20206020", -- 2f04
		x"00000000", -- 2f08
		x"00000000", -- 2f0c
		x"00000438", -- 2f10
		x"68282828", -- 2f14
		x"00000000", -- 2f18
		x"00000000", -- 2f1c
		x"f0f0f0f0", -- 2f20
		x"f0f0f0f0", -- 2f24
		x"f0f0f0f0", -- 2f28
		x"00000000", -- 2f2c
		x"0f0f0f0f", -- 2f30
		x"0f0f0f0f", -- 2f34
		x"0f0f0f0f", -- 2f38
		x"00000000", -- 2f3c
		x"ff818181", -- 2f40
		x"81818181", -- 2f44
		x"818181ff", -- 2f48
		x"00000000", -- 2f4c
		x"ffffffdf", -- 2f50
		x"bf00bfdf", -- 2f54
		x"ffffffff", -- 2f58
		x"00000000", -- 2f5c
		x"ffffff7f", -- 2f60
		x"bf1fbf7f", -- 2f64
		x"ffffffff", -- 2f68
		x"00000000", -- 2f6c
		x"fbf1eafb", -- 2f70
		x"fbfbfbfb", -- 2f74
		x"eaf1fbff", -- 2f78
		x"00000000", -- 2f7c
		x"ffffffff", -- 2f80
		x"83ffffff", -- 2f84
		x"ffffffff", -- 2f88
		x"00000000", -- 2f8c
		x"ffc7bbfb", -- 2f90
		x"f7efefff", -- 2f94
		x"efffffff", -- 2f98
		x"00000000", -- 2f9c
		x"ff1fbfbf", -- 2fa0
		x"bf19f6f6", -- 2fa4
		x"f6f9ffff", -- 2fa8
		x"00000000", -- 2fac
		x"ffffffff", -- 2fb0
		x"ffffffff", -- 2fb4
		x"ffffffff", -- 2fb8
		x"00000000", -- 2fbc
		x"00081838", -- 2fc0
		x"78381808", -- 2fc4
		x"00000000", -- 2fc8
		x"00000000", -- 2fcc
		x"ffffd7ef", -- 2fd0
		x"83efd7ff", -- 2fd4
		x"ffffffff", -- 2fd8
		x"00000000", -- 2fdc
		x"ff838383", -- 2fe0
		x"83838383", -- 2fe4
		x"ffffffff", -- 2fe8
		x"00000000", -- 2fec
		x"7cfebab6", -- 2ff0
		x"ae8eb6ba", -- 2ff4
		x"fe7c0000", -- 2ff8
		x"00000000", -- 2ffc
		x"00010203", -- 3000
		x"04050607", -- 3004
		x"08091011", -- 3008
		x"12131415", -- 300c
		x"16171819", -- 3010
		x"20212223", -- 3014
		x"24252627", -- 3018
		x"28293031", -- 301c
		x"32333435", -- 3020
		x"36373839", -- 3024
		x"40414243", -- 3028
		x"44454647", -- 302c
		x"48495051", -- 3030
		x"52535455", -- 3034
		x"56575859", -- 3038
		x"60616263", -- 303c
		x"64656667", -- 3040
		x"68697071", -- 3044
		x"72737475", -- 3048
		x"76777879", -- 304c
		x"80818283", -- 3050
		x"84858687", -- 3054
		x"88899091", -- 3058
		x"92939495", -- 305c
		x"96979899", -- 3060
		x"00010203", -- 3064
		x"04050607", -- 3068
		x"08090000", -- 306c
		x"00000001", -- 3070
		x"0a0b0c0d", -- 3074
		x"0e0f1011", -- 3078
		x"12130000", -- 307c
		x"00000000", -- 3080
		x"14151617", -- 3084
		x"18191a1b", -- 3088
		x"1c1d0000", -- 308c
		x"00000000", -- 3090
		x"1e1f2021", -- 3094
		x"22232425", -- 3098
		x"26270000", -- 309c
		x"00000000", -- 30a0
		x"28292a2b", -- 30a4
		x"2c2d2e2f", -- 30a8
		x"30310000", -- 30ac
		x"00000000", -- 30b0
		x"32333435", -- 30b4
		x"36373839", -- 30b8
		x"3a3b0000", -- 30bc
		x"00000000", -- 30c0
		x"3c3d3e3f", -- 30c4
		x"40414243", -- 30c8
		x"44450000", -- 30cc
		x"00000000", -- 30d0
		x"46474849", -- 30d4
		x"4a4b4c4d", -- 30d8
		x"4e4f0000", -- 30dc
		x"00000000", -- 30e0
		x"50515253", -- 30e4
		x"54555657", -- 30e8
		x"58590000", -- 30ec
		x"00000000", -- 30f0
		x"5a5b5c5d", -- 30f4
		x"5e5f6061", -- 30f8
		x"6263245f", -- 30fc
		x"201f205f", -- 3100
		x"225f2f0a", -- 3104
		x"4a806f42", -- 3108
		x"32083409", -- 310c
		x"02010001", -- 3110
		x"02020001", -- 3114
		x"b5016708", -- 3118
		x"10d95380", -- 311c
		x"6efa602a", -- 3120
		x"4a026706", -- 3124
		x"10d95380", -- 3128
		x"6f202200", -- 312c
		x"e4896706", -- 3130
		x"20d95381", -- 3134
		x"6efa0200", -- 3138
		x"00031200", -- 313c
		x"e2096702", -- 3140
		x"30d90200", -- 3144
		x"00016702", -- 3148
		x"10d94e75", -- 314c
		x"245f201f", -- 3150
		x"205f225f", -- 3154
		x"2f0a4a80", -- 3158
		x"6f46d1c0", -- 315c
		x"d3c03208", -- 3160
		x"34090201", -- 3164
		x"00010202", -- 3168
		x"0001b501", -- 316c
		x"67081121", -- 3170
		x"53806efa", -- 3174
		x"602a4a02", -- 3178
		x"67061121", -- 317c
		x"53806f20", -- 3180
		x"2200e489", -- 3184
		x"67062121", -- 3188
		x"53816efa", -- 318c
		x"02000003", -- 3190
		x"1200e209", -- 3194
		x"67023121", -- 3198
		x"02000001", -- 319c
		x"67021121", -- 31a0
		x"4e754cdf", -- 31a4
		x"00073041", -- 31a8
		x"b1c1660e", -- 31ac
		x"3042b1c2", -- 31b0
		x"6610c5c1", -- 31b4
		x"2f022040", -- 31b8
		x"4ed03042", -- 31bc
		x"b1c26634", -- 31c0
		x"c3423602", -- 31c4
		x"c6c12802", -- 31c8
		x"4844c8c1", -- 31cc
		x"48437a00", -- 31d0
		x"3a03d885", -- 31d4
		x"4a416a02", -- 31d8
		x"98824a82", -- 31dc
		x"6a063a01", -- 31e0
		x"48459885", -- 31e4
		x"3044b1c4", -- 31e8
		x"664e4843", -- 31ec
		x"3f033f04", -- 31f0
		x"20404ed0", -- 31f4
		x"26017e00", -- 31f8
		x"e2836402", -- 31fc
		x"2e023043", -- 3200
		x"b6886700", -- 3204
		x"00162602", -- 3208
		x"7e00e283", -- 320c
		x"64022e01", -- 3210
		x"3043b688", -- 3214
		x"66000022", -- 3218
		x"240143fa", -- 321c
		x"0008c189", -- 3220
		x"2203609e", -- 3224
		x"584fd643", -- 3228
		x"d984d647", -- 322c
		x"484748c7", -- 3230
		x"d9874843", -- 3234
		x"200960ac", -- 3238
		x"4e447e01", -- 323c
		x"60027e00", -- 3240
		x"4cdf0007", -- 3244
		x"4a81671a", -- 3248
		x"3041b288", -- 324c
		x"66162602", -- 3250
		x"87c16910", -- 3254
		x"4a476702", -- 3258
		x"484348c3", -- 325c
		x"2f032040", -- 3260
		x"4ed04e45", -- 3264
		x"780f7c00", -- 3268
		x"7a004a81", -- 326c
		x"6a064481", -- 3270
		x"69484646", -- 3274
		x"4a826a10", -- 3278
		x"44826808", -- 327c
		x"b2bcffff", -- 3280
		x"ffff67b4", -- 3284
		x"46464645", -- 3288
		x"76004841", -- 328c
		x"4a41663c", -- 3290
		x"48424841", -- 3294
		x"360286c1", -- 3298
		x"34034842", -- 329c
		x"360286c1", -- 32a0
		x"34034243", -- 32a4
		x"48434a46", -- 32a8
		x"6a024482", -- 32ac
		x"4a456a02", -- 32b0
		x"44834a47", -- 32b4
		x"66a6c543", -- 32b8
		x"60a24482", -- 32bc
		x"69082602", -- 32c0
		x"44837400", -- 32c4
		x"60ec7401", -- 32c8
		x"760060e6", -- 32cc
		x"48414842", -- 32d0
		x"36024242", -- 32d4
		x"96812041", -- 32d8
		x"4481d482", -- 32dc
		x"d783d688", -- 32e0
		x"6a1251cc", -- 32e4
		x"fff6d688", -- 32e8
		x"d48260ba", -- 32ec
		x"d582d783", -- 32f0
		x"d6816bee", -- 32f4
		x"51ccfff6", -- 32f8
		x"d58260aa", -- 32fc
		x"1f3c0001", -- 3300
		x"1f3c0000", -- 3304
		x"60081f3c", -- 3308
		x"00001f3c", -- 330c
		x"0001266f", -- 3310
		x"0008286f", -- 3314
		x"000c3e1b", -- 3318
		x"3c1cbe46", -- 331c
		x"6f043a06", -- 3320
		x"60023a07", -- 3324
		x"6714e445", -- 3328
		x"6408b94b", -- 332c
		x"662c4a45", -- 3330
		x"6708b98b", -- 3334
		x"66245345", -- 3338
		x"6ef89e46", -- 333c
		x"67166a0c", -- 3340
		x"44474a5c", -- 3344
		x"66145547", -- 3348
		x"6ef86008", -- 334c
		x"4a5b660a", -- 3350
		x"55476ef8", -- 3354
		x"1f57000e", -- 3358
		x"60061f6f", -- 335c
		x"0002000e", -- 3360
		x"2f6f0004", -- 3364
		x"000adffc", -- 3368
		x"0000000a", -- 336c
		x"4e75266f", -- 3370
		x"0004286f", -- 3374
		x"00083e1b", -- 3378
		x"38c76710", -- 337c
		x"e4476406", -- 3380
		x"38db4a47", -- 3384
		x"670628db", -- 3388
		x"53476efa", -- 338c
		x"2f570008", -- 3390
		x"508f4e75", -- 3394
		x"246f0004", -- 3398
		x"286f0008", -- 339c
		x"266f000c", -- 33a0
		x"3e1a3c1c", -- 33a4
		x"be466f06", -- 33a8
		x"3a0636c7", -- 33ac
		x"60043a07", -- 33b0
		x"36c64a45", -- 33b4
		x"6718e445", -- 33b8
		x"640a381a", -- 33bc
		x"885c36c4", -- 33c0
		x"4a45670a", -- 33c4
		x"281a889c", -- 33c8
		x"26c45345", -- 33cc
		x"6ef69e46", -- 33d0
		x"67126a0a", -- 33d4
		x"444736dc", -- 33d8
		x"55476efa", -- 33dc
		x"600636da", -- 33e0
		x"55476efa", -- 33e4
		x"2f57000c", -- 33e8
		x"dffc0000", -- 33ec
		x"000c4e75", -- 33f0
		x"266f0004", -- 33f4
		x"286f0008", -- 33f8
		x"3e1b3c1c", -- 33fc
		x"be466f04", -- 3400
		x"3a066002", -- 3404
		x"3a07671c", -- 3408
		x"e445640c", -- 340c
		x"381b4644", -- 3410
		x"c85c6624", -- 3414
		x"4a45670c", -- 3418
		x"281b4684", -- 341c
		x"c89c6618", -- 3420
		x"53456ef4", -- 3424
		x"9c476f08", -- 3428
		x"4a5c660c", -- 342c
		x"55466ef8", -- 3430
		x"1f7c0001", -- 3434
		x"000a6006", -- 3438
		x"1f7c0000", -- 343c
		x"000a2f57", -- 3440
		x"00065c8f", -- 3444
		x"4e75246f", -- 3448
		x"0004286f", -- 344c
		x"0008266f", -- 3450
		x"000c3e1a", -- 3454
		x"be5c6f04", -- 3458
		x"3e2cfffe", -- 345c
		x"36c76718", -- 3460
		x"e447640a", -- 3464
		x"3c1acc5c", -- 3468
		x"36c64a47", -- 346c
		x"670a2c1a", -- 3470
		x"cc9c26c6", -- 3474
		x"53476ef6", -- 3478
		x"2f57000c", -- 347c
		x"dffc0000", -- 3480
		x"000c4e75", -- 3484
		x"246f0004", -- 3488
		x"286f0008", -- 348c
		x"266f000c", -- 3490
		x"3e1a3c1c", -- 3494
		x"be466f04", -- 3498
		x"3a066002", -- 349c
		x"3a0736c6", -- 34a0
		x"4a45671c", -- 34a4
		x"e445640c", -- 34a8
		x"381a4644", -- 34ac
		x"c85c36c4", -- 34b0
		x"4a45670c", -- 34b4
		x"281a4684", -- 34b8
		x"c89c26c4", -- 34bc
		x"53456ef4", -- 34c0
		x"9c476f06", -- 34c4
		x"36dc5546", -- 34c8
		x"6efa2f57", -- 34cc
		x"000cdffc", -- 34d0
		x"0000000c", -- 34d4
		x"4e75205f", -- 34d8
		x"225f201f", -- 34dc
		x"6d1881fc", -- 34e0
		x"0008b051", -- 34e4
		x"6c102200", -- 34e8
		x"48411031", -- 34ec
		x"0002e328", -- 34f0
		x"ee081f00", -- 34f4
		x"4ed04227", -- 34f8
		x"4ed0205f", -- 34fc
		x"301f225f", -- 3500
		x"24573e19", -- 3504
		x"34c7b3ca", -- 3508
		x"670c264a", -- 350c
		x"3c076f06", -- 3510
		x"36d95546", -- 3514
		x"6efa48c0", -- 3518
		x"81fc0010", -- 351c
		x"2a004845", -- 3520
		x"9a7c000f", -- 3524
		x"4445e340", -- 3528
		x"32005441", -- 352c
		x"3401926a", -- 3530
		x"fffe6f0e", -- 3534
		x"3542fffe", -- 3538
		x"47f22000", -- 353c
		x"42635541", -- 3540
		x"6efa0885", -- 3544
		x"00036706", -- 3548
		x"0bf20000", -- 354c
		x"4ed00bf2", -- 3550
		x"00014ed0", -- 3554
		x"4cdf1c00", -- 3558
		x"4244181b", -- 355c
		x"67164245", -- 3560
		x"1a1443f4", -- 3564
		x"5001da04", -- 3568
		x"650a1885", -- 356c
		x"534412db", -- 3570
		x"51ccfffc", -- 3574
		x"4ed2245f", -- 3578
		x"2e1f285f", -- 357c
		x"265f6f32", -- 3580
		x"4244181b", -- 3584
		x"672c4245", -- 3588
		x"1a1443f4", -- 358c
		x"50013605", -- 3590
		x"da04651e", -- 3594
		x"18859647", -- 3598
		x"6c065243", -- 359c
		x"670e4ed2", -- 35a0
		x"41f14000", -- 35a4
		x"112151cb", -- 35a8
		x"fffc5344", -- 35ac
		x"12db51cc", -- 35b0
		x"fffc4ed2", -- 35b4
		x"245f2c1f", -- 35b8
		x"2e1f265f", -- 35bc
		x"285f6f24", -- 35c0
		x"4a866d20", -- 35c4
		x"42441813", -- 35c8
		x"52449847", -- 35cc
		x"6d16bc44", -- 35d0
		x"6f023c04", -- 35d4
		x"18c65346", -- 35d8
		x"6d0a43f3", -- 35dc
		x"700018d9", -- 35e0
		x"51cefffc", -- 35e4
		x"4ed2245f", -- 35e8
		x"2c1f2e1f", -- 35ec
		x"285f6f28", -- 35f0
		x"4a866f24", -- 35f4
		x"42451a14", -- 35f8
		x"9a466d1c", -- 35fc
		x"36055243", -- 3600
		x"96476d14", -- 3604
		x"18855343", -- 3608
		x"6d0e43f4", -- 360c
		x"700041f1", -- 3610
		x"600012d8", -- 3614
		x"51cbfffc", -- 3618
		x"4ed24cdf", -- 361c
		x"1c004297", -- 3620
		x"42451a1c", -- 3624
		x"672c4284", -- 3628
		x"181b9845", -- 362c
		x"6d24101c", -- 3630
		x"55452204", -- 3634
		x"b01b57cc", -- 3638
		x"fffc6616", -- 363c
		x"34056d0c", -- 3640
		x"43d441d3", -- 3644
		x"b10956ca", -- 3648
		x"fffc66ea", -- 364c
		x"92445241", -- 3650
		x"2e814ed2", -- 3654
		x"2f52f8ac", -- 3658
		x"174d6123", -- 365c
		x"2f87b6d7", -- 3660
		x"1d20b96c", -- 3664
		x"2fbda48c", -- 3668
		x"e468e7c7", -- 366c
		x"2ff286d8", -- 3670
		x"0ec190dc", -- 3674
		x"3027288e", -- 3678
		x"1271f513", -- 367c
		x"305cf2b1", -- 3680
		x"970e7258", -- 3684
		x"309217ae", -- 3688
		x"fe690777", -- 368c
		x"30c69d9a", -- 3690
		x"be034955", -- 3694
		x"30fc4501", -- 3698
		x"6d841baa", -- 369c
		x"3131ab20", -- 36a0
		x"e472914a", -- 36a4
		x"316615e9", -- 36a8
		x"1d8f359d", -- 36ac
		x"319b9b63", -- 36b0
		x"64f30304", -- 36b4
		x"31d1411e", -- 36b8
		x"1f17e1e3", -- 36bc
		x"32059165", -- 36c0
		x"a6ddda5b", -- 36c4
		x"323af5bf", -- 36c8
		x"109550f2", -- 36cc
		x"3270d997", -- 36d0
		x"6a5d5297", -- 36d4
		x"32a50ffd", -- 36d8
		x"44f4a73d", -- 36dc
		x"32da53fc", -- 36e0
		x"9631d10d", -- 36e4
		x"3310747d", -- 36e8
		x"dddf22a8", -- 36ec
		x"3344919d", -- 36f0
		x"5556eb52", -- 36f4
		x"3379b604", -- 36f8
		x"aaaca626", -- 36fc
		x"33b011c2", -- 3700
		x"eaabe7d8", -- 3704
		x"33e41633", -- 3708
		x"a556e1ce", -- 370c
		x"34191bc0", -- 3710
		x"8eac9a41", -- 3714
		x"344f62b0", -- 3718
		x"b257c0d2", -- 371c
		x"34839dae", -- 3720
		x"6f76d883", -- 3724
		x"34b8851a", -- 3728
		x"0b548ea4", -- 372c
		x"34eea660", -- 3730
		x"8e29b24d", -- 3734
		x"352327fc", -- 3738
		x"58da0f70", -- 373c
		x"3557f1fb", -- 3740
		x"6f10934c", -- 3744
		x"358dee7a", -- 3748
		x"4ad4b81f", -- 374c
		x"35c2b50c", -- 3750
		x"6ec4f313", -- 3754
		x"35f7624f", -- 3758
		x"8a762fd8", -- 375c
		x"362d3ae3", -- 3760
		x"6d13bbce", -- 3764
		x"366244ce", -- 3768
		x"242c5561", -- 376c
		x"3696d601", -- 3770
		x"ad376ab9", -- 3774
		x"36cc8b82", -- 3778
		x"18854567", -- 377c
		x"3701d731", -- 3780
		x"4f534b61", -- 3784
		x"37364cfd", -- 3788
		x"a3281e39", -- 378c
		x"376be03d", -- 3790
		x"0bf225c7", -- 3794
		x"37a16c26", -- 3798
		x"2777579c", -- 379c
		x"37d5c72f", -- 37a0
		x"b1552d83", -- 37a4
		x"380b38fb", -- 37a8
		x"9daa78e4", -- 37ac
		x"3841039d", -- 37b0
		x"428a8b8f", -- 37b4
		x"38754484", -- 37b8
		x"932d2e72", -- 37bc
		x"38aa95a5", -- 37c0
		x"b7f87a0f", -- 37c4
		x"38e09d87", -- 37c8
		x"92fb4c49", -- 37cc
		x"3914c4e9", -- 37d0
		x"77ba1f5c", -- 37d4
		x"3949f623", -- 37d8
		x"d5a8a733", -- 37dc
		x"398039d6", -- 37e0
		x"65896880", -- 37e4
		x"39b4484b", -- 37e8
		x"feebc2a0", -- 37ec
		x"39e95a5e", -- 37f0
		x"fea6b347", -- 37f4
		x"3a1fb0f6", -- 37f8
		x"be506019", -- 37fc
		x"3a53ce9a", -- 3800
		x"36f23c10", -- 3804
		x"3a88c240", -- 3808
		x"c4aecb14", -- 380c
		x"3abef2d0", -- 3810
		x"f5da7dd9", -- 3814
		x"3af357c2", -- 3818
		x"99a88ea7", -- 381c
		x"3b282db3", -- 3820
		x"4012b251", -- 3824
		x"3b5e3920", -- 3828
		x"10175ee6", -- 382c
		x"3b92e3b4", -- 3830
		x"0a0e9b4f", -- 3834
		x"3bc79ca1", -- 3838
		x"0c924223", -- 383c
		x"3bfd83c9", -- 3840
		x"4fb6d2ac", -- 3844
		x"3c32725d", -- 3848
		x"d1d243ac", -- 384c
		x"3c670ef5", -- 3850
		x"4646d497", -- 3854
		x"3c9cd2b2", -- 3858
		x"97d889bc", -- 385c
		x"3cd203af", -- 3860
		x"9ee75616", -- 3864
		x"3d06849b", -- 3868
		x"86a12b9b", -- 386c
		x"3d3c25c2", -- 3870
		x"68497682", -- 3874
		x"3d719799", -- 3878
		x"812dea11", -- 387c
		x"3da5fd7f", -- 3880
		x"e1796495", -- 3884
		x"3ddb7cdf", -- 3888
		x"d9d7bdbb", -- 388c
		x"3e112e0b", -- 3890
		x"e826d695", -- 3894
		x"3e45798e", -- 3898
		x"e2308c3a", -- 389c
		x"3e7ad7f2", -- 38a0
		x"9abcaf48", -- 38a4
		x"3eb0c6f7", -- 38a8
		x"a0b5ed8d", -- 38ac
		x"3ee4f8b5", -- 38b0
		x"88e368f1", -- 38b4
		x"3f1a36e2", -- 38b8
		x"eb1c432d", -- 38bc
		x"3f50624d", -- 38c0
		x"d2f1a9fc", -- 38c4
		x"3f847ae1", -- 38c8
		x"47ae147b", -- 38cc
		x"3fb99999", -- 38d0
		x"9999999a", -- 38d4
		x"3ff00000", -- 38d8
		x"00000000", -- 38dc
		x"40240000", -- 38e0
		x"00000000", -- 38e4
		x"40590000", -- 38e8
		x"00000000", -- 38ec
		x"408f4000", -- 38f0
		x"00000000", -- 38f4
		x"40c38800", -- 38f8
		x"00000000", -- 38fc
		x"40f86a00", -- 3900
		x"00000000", -- 3904
		x"412e8480", -- 3908
		x"00000000", -- 390c
		x"416312d0", -- 3910
		x"00000000", -- 3914
		x"4197d784", -- 3918
		x"00000000", -- 391c
		x"41cdcd65", -- 3920
		x"00000000", -- 3924
		x"4202a05f", -- 3928
		x"20000000", -- 392c
		x"42374876", -- 3930
		x"e8000000", -- 3934
		x"426d1a94", -- 3938
		x"a2000000", -- 393c
		x"42a2309c", -- 3940
		x"e5400000", -- 3944
		x"42d6bcc4", -- 3948
		x"1e900000", -- 394c
		x"430c6bf5", -- 3950
		x"26340000", -- 3954
		x"4341c379", -- 3958
		x"37e08000", -- 395c
		x"43763457", -- 3960
		x"85d8a000", -- 3964
		x"43abc16d", -- 3968
		x"674ec800", -- 396c
		x"43e158e4", -- 3970
		x"60913d00", -- 3974
		x"4415af1d", -- 3978
		x"78b58c40", -- 397c
		x"444b1ae4", -- 3980
		x"d6e2ef50", -- 3984
		x"4480f0cf", -- 3988
		x"064dd592", -- 398c
		x"44b52d02", -- 3990
		x"c7e14af6", -- 3994
		x"44ea7843", -- 3998
		x"79d99db4", -- 399c
		x"45208b2a", -- 39a0
		x"2c280291", -- 39a4
		x"4554adf4", -- 39a8
		x"b7320335", -- 39ac
		x"4589d971", -- 39b0
		x"e4fe8402", -- 39b4
		x"45c027e7", -- 39b8
		x"2f1f1281", -- 39bc
		x"45f431e0", -- 39c0
		x"fae6d721", -- 39c4
		x"46293e59", -- 39c8
		x"39a08cea", -- 39cc
		x"465f8def", -- 39d0
		x"8808b024", -- 39d4
		x"4693b8b5", -- 39d8
		x"b5056e17", -- 39dc
		x"46c8a6e3", -- 39e0
		x"2246c99c", -- 39e4
		x"46fed09b", -- 39e8
		x"ead87c03", -- 39ec
		x"47334261", -- 39f0
		x"72c74d82", -- 39f4
		x"476812f9", -- 39f8
		x"cf7920e3", -- 39fc
		x"479e17b8", -- 3a00
		x"4357691b", -- 3a04
		x"47d2ced3", -- 3a08
		x"2a16a1b1", -- 3a0c
		x"48078287", -- 3a10
		x"f49c4a1d", -- 3a14
		x"483d6329", -- 3a18
		x"f1c35ca5", -- 3a1c
		x"48725dfa", -- 3a20
		x"371a19e7", -- 3a24
		x"48a6f578", -- 3a28
		x"c4e0a061", -- 3a2c
		x"48dcb2d6", -- 3a30
		x"f618c879", -- 3a34
		x"4911efc6", -- 3a38
		x"59cf7d4c", -- 3a3c
		x"49466bb7", -- 3a40
		x"f0435c9e", -- 3a44
		x"497c06a5", -- 3a48
		x"ec5433c6", -- 3a4c
		x"49b18427", -- 3a50
		x"b3b4a05c", -- 3a54
		x"49e5e531", -- 3a58
		x"a0a1c873", -- 3a5c
		x"4a1b5e7e", -- 3a60
		x"08ca3a8f", -- 3a64
		x"4a511b0e", -- 3a68
		x"c57e649a", -- 3a6c
		x"4a8561d2", -- 3a70
		x"76ddfdc0", -- 3a74
		x"4ababa47", -- 3a78
		x"14957d30", -- 3a7c
		x"4af0b46c", -- 3a80
		x"6cdd6e3e", -- 3a84
		x"4b24e187", -- 3a88
		x"8814c9ce", -- 3a8c
		x"4b5a19e9", -- 3a90
		x"6a19fc41", -- 3a94
		x"4b905031", -- 3a98
		x"e2503da9", -- 3a9c
		x"4bc4643e", -- 3aa0
		x"5ae44d13", -- 3aa4
		x"4bf97d4d", -- 3aa8
		x"f19d6057", -- 3aac
		x"4c2fdca1", -- 3ab0
		x"6e04b86d", -- 3ab4
		x"4c63e9e4", -- 3ab8
		x"e4c2f344", -- 3abc
		x"4c98e45e", -- 3ac0
		x"1df3b015", -- 3ac4
		x"4ccf1d75", -- 3ac8
		x"a5709c1b", -- 3acc
		x"4d037269", -- 3ad0
		x"87666191", -- 3ad4
		x"4d384f03", -- 3ad8
		x"e93ff9f5", -- 3adc
		x"0ac80628", -- 3ae0
		x"64ac6f43", -- 3ae4
		x"18123ff0", -- 3ae8
		x"6eea847a", -- 3aec
		x"255bba08", -- 3af0
		x"cf8c979d", -- 3af4
		x"32a50ffd", -- 3af8
		x"44f4a73d", -- 3afc
		x"3ff00000", -- 3b00
		x"00000000", -- 3b04
		x"4d384f03", -- 3b08
		x"e93ff9f5", -- 3b0c
		x"5a827748", -- 3b10
		x"f9301d32", -- 3b14
		x"67cc0e1e", -- 3b18
		x"f1a724eb", -- 3b1c
		x"75154fdd", -- 3b20
		x"7f73bf3c", -- 3b24
		x"00010203", -- 3b28
		x"04050607", -- 3b2c
		x"08090000", -- 3b30
		x"00000000", -- 3b34
		x"0a0b0c0d", -- 3b38
		x"0e0f1011", -- 3b3c
		x"12130000", -- 3b40
		x"00000000", -- 3b44
		x"14151617", -- 3b48
		x"18191a1b", -- 3b4c
		x"1c1d0000", -- 3b50
		x"00000000", -- 3b54
		x"1e1f2021", -- 3b58
		x"22232425", -- 3b5c
		x"26270000", -- 3b60
		x"00000000", -- 3b64
		x"28292a2b", -- 3b68
		x"2c2d2e2f", -- 3b6c
		x"30310000", -- 3b70
		x"00000000", -- 3b74
		x"32333435", -- 3b78
		x"36373839", -- 3b7c
		x"3a3b0000", -- 3b80
		x"00000000", -- 3b84
		x"3c3d3e3f", -- 3b88
		x"40414243", -- 3b8c
		x"44450000", -- 3b90
		x"00000000", -- 3b94
		x"46474849", -- 3b98
		x"4a4b4c4d", -- 3b9c
		x"4e4f0000", -- 3ba0
		x"00000000", -- 3ba4
		x"50515253", -- 3ba8
		x"54555657", -- 3bac
		x"58590000", -- 3bb0
		x"00000000", -- 3bb4
		x"5a5b5c5d", -- 3bb8
		x"5e5f6061", -- 3bbc
		x"62630001", -- 3bc0
		x"02030405", -- 3bc4
		x"06070809", -- 3bc8
		x"10111213", -- 3bcc
		x"14151617", -- 3bd0
		x"18192021", -- 3bd4
		x"22232425", -- 3bd8
		x"26272829", -- 3bdc
		x"30313233", -- 3be0
		x"34353637", -- 3be4
		x"38394041", -- 3be8
		x"42434445", -- 3bec
		x"46474849", -- 3bf0
		x"50515253", -- 3bf4
		x"54555657", -- 3bf8
		x"58596061", -- 3bfc
		x"62636465", -- 3c00
		x"66676869", -- 3c04
		x"70717273", -- 3c08
		x"74757677", -- 3c0c
		x"78798081", -- 3c10
		x"82838485", -- 3c14
		x"86878889", -- 3c18
		x"90919293", -- 3c1c
		x"94959697", -- 3c20
		x"9899bfe9", -- 3c24
		x"4415b356", -- 3c28
		x"bd294030", -- 3c2c
		x"624a2016", -- 3c30
		x"afedc050", -- 3c34
		x"07ff12b3", -- 3c38
		x"b59ac041", -- 3c3c
		x"d5804b67", -- 3c40
		x"ce0f4073", -- 3c44
		x"8083fa15", -- 3c48
		x"267ec088", -- 3c4c
		x"0bfe9c0d", -- 3c50
		x"90773f00", -- 3c54
		x"8b442ae6", -- 3c58
		x"921e3f7f", -- 3c5c
		x"074bf22a", -- 3c60
		x"12a63fd0", -- 3c64
		x"00000000", -- 3c68
		x"00003ea9", -- 3c6c
		x"33630ce5", -- 3c70
		x"04553f44", -- 3c74
		x"af0c5c28", -- 3c78
		x"d4df3fad", -- 3c7c
		x"172851df", -- 3c80
		x"d9ff3fe0", -- 3c84
		x"00000000", -- 3c88
		x"00003ce8", -- 3c8c
		x"80ff6993", -- 3c90
		x"df95bd6a", -- 3c94
		x"e420dc08", -- 3c98
		x"499c3de6", -- 3c9c
		x"123c686a", -- 3ca0
		x"d430be5a", -- 3ca4
		x"e6454b5d", -- 3ca8
		x"c0ab3ec7", -- 3cac
		x"1de3a524", -- 3cb0
		x"f063bf2a", -- 3cb4
		x"01a01a01", -- 3cb8
		x"3e1a3f81", -- 3cbc
		x"11111111", -- 3cc0
		x"10b0bfc5", -- 3cc4
		x"55555555", -- 3cc8
		x"5555bef2", -- 3ccc
		x"bab72ea2", -- 3cd0
		x"c7243f6c", -- 3cd4
		x"0e82a63b", -- 3cd8
		x"aadfbfc1", -- 3cdc
		x"12b5e54d", -- 3ce0
		x"09003ff0", -- 3ce4
		x"00000000", -- 3ce8
		x"00003ea0", -- 3cec
		x"b774f076", -- 3cf0
		x"78e9bf34", -- 3cf4
		x"6f649909", -- 3cf8
		x"48413f9a", -- 3cfc
		x"479ea17e", -- 3d00
		x"2159bfdd", -- 3d04
		x"deb047fb", -- 3d08
		x"d9d53ff0", -- 3d0c
		x"00000000", -- 3d10
		x"0000bfe6", -- 3d14
		x"4bbdb5e6", -- 3d18
		x"1e654024", -- 3d1c
		x"4e1764ec", -- 3d20
		x"3927c043", -- 3d24
		x"d82ca9a6", -- 3d28
		x"da9f404c", -- 3d2c
		x"9aa7360a", -- 3d30
		x"d48ac03b", -- 3d34
		x"5e55a83a", -- 3d38
		x"0a62c037", -- 3d3c
		x"d2e86ef9", -- 3d40
		x"861f4062", -- 3d44
		x"de7c9659", -- 3d48
		x"1c70c077", -- 3d4c
		x"ddcefc56", -- 3d50
		x"a848407a", -- 3d54
		x"124f101e", -- 3d58
		x"b843c064", -- 3d5c
		x"86c03e2b", -- 3d60
		x"87ccbfea", -- 3d64
		x"cd7ad9b1", -- 3d68
		x"87bdc020", -- 3d6c
		x"fd3f5c8d", -- 3d70
		x"6a63c034", -- 3d74
		x"817fb9e2", -- 3d78
		x"bccbc02b", -- 3d7c
		x"60a65106", -- 3d80
		x"1ce2402e", -- 3d84
		x"0c49e14a", -- 3d88
		x"c710404d", -- 3d8c
		x"ca0a320d", -- 3d90
		x"a3d74055", -- 3d94
		x"8a12040b", -- 3d98
		x"6da54044", -- 3d9c
		x"887cbcc4", -- 3da0
		x"95a93f3c", -- 3da4
		x"78fddb4a", -- 3da8
		x"fc283f62", -- 3dac
		x"49242e27", -- 3db0
		x"8dac3f89", -- 3db4
		x"9999999e", -- 3db8
		x"080e3fb5", -- 3dbc
		x"55555555", -- 3dc0
		x"554d3eef", -- 3dc4
		x"4edde392", -- 3dc8
		x"cc803f24", -- 3dcc
		x"2f7ae038", -- 3dd0
		x"4c743f55", -- 3dd4
		x"d87e18d7", -- 3dd8
		x"cd9f3f83", -- 3ddc
		x"b2ab6e13", -- 3de0
		x"1d983fac", -- 3de4
		x"6b08d703", -- 3de8
		x"026d3fce", -- 3dec
		x"bfbdff82", -- 3df0
		x"c4ce3fe6", -- 3df4
		x"2e42fefa", -- 3df8
		x"39ef0000", -- 3dfc
		x"00000000", -- 3e00
		x"00003ff0", -- 3e04
		x"00000000", -- 3e08
		x"00003fee", -- 3e0c
		x"a4afa2a4", -- 3e10
		x"90da3fed", -- 3e14
		x"5818dcfb", -- 3e18
		x"a4873fec", -- 3e1c
		x"199bdd85", -- 3e20
		x"529c3fea", -- 3e24
		x"e89f995a", -- 3e28
		x"d3ad3fe9", -- 3e2c
		x"c49182a3", -- 3e30
		x"f0903fe8", -- 3e34
		x"ace5422a", -- 3e38
		x"a0db3fe7", -- 3e3c
		x"a11473eb", -- 3e40
		x"01873fe6", -- 3e44
		x"a09e667f", -- 3e48
		x"3bcd3fe5", -- 3e4c
		x"ab07dd48", -- 3e50
		x"54293fe4", -- 3e54
		x"bfdad536", -- 3e58
		x"2a273fe3", -- 3e5c
		x"dea64c12", -- 3e60
		x"34223fe3", -- 3e64
		x"06fe0a31", -- 3e68
		x"b7153fe2", -- 3e6c
		x"387a6e75", -- 3e70
		x"62383fe1", -- 3e74
		x"72b83c7d", -- 3e78
		x"517b3fe0", -- 3e7c
		x"b5586cf9", -- 3e80
		x"890f3fe0", -- 3e84
		x"00000000", -- 3e88
		x"00000000", -- 3e8c
		x"00000000", -- 3e90
		x"0000bc7e", -- 3e94
		x"9c23179c", -- 3e98
		x"00003c61", -- 3e9c
		x"10658950", -- 3ea0
		x"00003c5c", -- 3ea4
		x"7c46b070", -- 3ea8
		x"0000bc64", -- 3eac
		x"1577ee04", -- 3eb0
		x"00003c76", -- 3eb4
		x"324c0546", -- 3eb8
		x"00003c6a", -- 3ebc
		x"da0911f0", -- 3ec0
		x"00003c79", -- 3ec4
		x"b07eb6c8", -- 3ec8
		x"00003c78", -- 3ecc
		x"a62e4adc", -- 3ed0
		x"00004e75", -- 3ed4
		x"2878fed4", -- 3ed8
		x"08380006", -- 3edc
		x"fed2665c", -- 3ee0
		x"08ac0000", -- 3ee4
		x"005c7000", -- 3ee8
		x"61000f46", -- 3eec
		x"4a6c00a0", -- 3ef0
		x"6b0c102c", -- 3ef4
		x"00a14640", -- 3ef8
		x"13c00001", -- 3efc
		x"ffff102c", -- 3f00
		x"00a10c00", -- 3f04
		x"000e6642", -- 3f08
		x"4a2c00a9", -- 3f0c
		x"670641fa", -- 3f10
		x"1af86004", -- 3f14
		x"41fa1ac8", -- 3f18
		x"610018ae", -- 3f1c
		x"08ec0002", -- 3f20
		x"005c08ac", -- 3f24
		x"0006000a", -- 3f28
		x"102c00a1", -- 3f2c
		x"6100109e", -- 3f30
		x"082c0002", -- 3f34
		x"005c66f8", -- 3f38
		x"6000008a", -- 3f3c
		x"08ec0000", -- 3f40
		x"005c08b8", -- 3f44
		x"0006fed2", -- 3f48
		x"609c082c", -- 3f4c
		x"0000005c", -- 3f50
		x"66724a2c", -- 3f54
		x"00a1676c", -- 3f58
		x"4a2c00a9", -- 3f5c
		x"670641fa", -- 3f60
		x"1afb6004", -- 3f64
		x"41fa1acd", -- 3f68
		x"6100185e", -- 3f6c
		x"4dfac966", -- 3f70
		x"08ec0002", -- 3f74
		x"005c08ac", -- 3f78
		x"0006000a", -- 3f7c
		x"102c00a1", -- 3f80
		x"6100104a", -- 3f84
		x"08380001", -- 3f88
		x"feda6620", -- 3f8c
		x"48790393", -- 3f90
		x"87004857", -- 3f94
		x"4eba1284", -- 3f98
		x"082c0002", -- 3f9c
		x"005c6708", -- 3fa0
		x"48574eba", -- 3fa4
		x"12966af0", -- 3fa8
		x"588f6012", -- 3fac
		x"223c008c", -- 3fb0
		x"d9d0082c", -- 3fb4
		x"0002005c", -- 3fb8
		x"67045381", -- 3fbc
		x"6ef408ac", -- 3fc0
		x"0002005c", -- 3fc4
		x"08ec0006", -- 3fc8
		x"000a4e75", -- 3fcc
		x"424f4f54", -- 3fd0
		x"524f4d20", -- 3fd4
		x"5265762e", -- 3fd8
		x"20440000", -- 3fdc
		x"ffffffff", -- 3fe0
		x"ffffffff", -- 3fe4
		x"ffffffff", -- 3fe8
		x"ffffffff", -- 3fec
		x"ffffffff", -- 3ff0
		x"f096a5c3", -- 3ff4
		x"db247a25", -- 3ff8
		x"0007000d", -- 3ffc
		x"4efa00fc", -- 4000
		x"4efa10f8", -- 4004
		x"4efa113c", -- 4008
		x"4efa115e", -- 400c
		x"4efa1182", -- 4010
		x"4efa10dc", -- 4014
		x"4efa10de", -- 4018
		x"7baa3e8d", -- 401c
		x"000051b8", -- 4020
		x"00000004", -- 4024
		x"0000474a", -- 4028
		x"00000004", -- 402c
		x"0000478c", -- 4030
		x"00000004", -- 4034
		x"000051c8", -- 4038
		x"00000004", -- 403c
		x"000045a4", -- 4040
		x"00000004", -- 4044
		x"000045c6", -- 4048
		x"00000004", -- 404c
		x"000051c0", -- 4050
		x"00000004", -- 4054
		x"00004752", -- 4058
		x"00000004", -- 405c
		x"00004794", -- 4060
		x"00000004", -- 4064
		x"000051d0", -- 4068
		x"00000004", -- 406c
		x"000045ac", -- 4070
		x"00000004", -- 4074
		x"00000000", -- 4078
		x"0000000a", -- 407c
		x"0000d4a4", -- 4080
		x"00000000", -- 4084
		x"000a0000", -- 4088
		x"d4a42000", -- 408c
		x"0000000a", -- 4090
		x"0000d4a4", -- 4094
		x"40000000", -- 4098
		x"000a0000", -- 409c
		x"45b4e000", -- 40a0
		x"0000000a", -- 40a4
		x"00004736", -- 40a8
		x"e1000000", -- 40ac
		x"000a0000", -- 40b0
		x"4778e200", -- 40b4
		x"00000000", -- 40b8
		x"00004478", -- 40bc
		x"000031fc", -- 40c0
		x"000cfdc0", -- 40c4
		x"4a38fdc2", -- 40c8
		x"672008f8", -- 40cc
		x"0002fdcc", -- 40d0
		x"4a38fdc3", -- 40d4
		x"6600c674", -- 40d8
		x"08b80002", -- 40dc
		x"fdcc21fc", -- 40e0
		x"e0ffffff", -- 40e4
		x"fedc6000", -- 40e8
		x"c6624278", -- 40ec
		x"fdc06000", -- 40f0
		x"c65a31fc", -- 40f4
		x"0012fdc0", -- 40f8
		x"60ca48e7", -- 40fc
		x"87984e55", -- 4100
		x"ffe82f38", -- 4104
		x"fffc6100", -- 4108
		x"09e821fc", -- 410c
		x"000043a4", -- 4110
		x"fffc487a", -- 4114
		x"02522b4f", -- 4118
		x"fff62878", -- 411c
		x"fed4302c", -- 4120
		x"00565340", -- 4124
		x"610015f0", -- 4128
		x"41fa17d0", -- 412c
		x"610015c6", -- 4130
		x"48e7fff8", -- 4134
		x"558f2f2d", -- 4138
		x"00286100", -- 413c
		x"2db66100", -- 4140
		x"0fba6100", -- 4144
		x"2dc24a1f", -- 4148
		x"4cdf1fff", -- 414c
		x"67000200", -- 4150
		x"48e7fff8", -- 4154
		x"558f2f2d", -- 4158
		x"0024486d", -- 415c
		x"fff2486d", -- 4160
		x"ffee3b7c", -- 4164
		x"e942ffe8", -- 4168
		x"486dffe8", -- 416c
		x"61002d84", -- 4170
		x"61000fd0", -- 4174
		x"61002d90", -- 4178
		x"4a1f4cdf", -- 417c
		x"1fff6700", -- 4180
		x"01ce4aad", -- 4184
		x"ffee6700", -- 4188
		x"00b04285", -- 418c
		x"420748e7", -- 4190
		x"fff82f05", -- 4194
		x"48780100", -- 4198
		x"4878fdd2", -- 419c
		x"42276100", -- 41a0
		x"2d526100", -- 41a4
		x"0fc46100", -- 41a8
		x"2d5e4cdf", -- 41ac
		x"1fff2678", -- 41b0
		x"fdd22c38", -- 41b4
		x"fdd62006", -- 41b8
		x"204bd088", -- 41bc
		x"650001da", -- 41c0
		x"b0bcffff", -- 41c4
		x"fac06200", -- 41c8
		x"01d0b0b8", -- 41cc
		x"fed46308", -- 41d0
		x"b7f8fdce", -- 41d4
		x"650001ca", -- 41d8
		x"50c75285", -- 41dc
		x"41f8fdda", -- 41e0
		x"bcbc0000", -- 41e4
		x"00f86e0a", -- 41e8
		x"4a866f3e", -- 41ec
		x"16d85386", -- 41f0
		x"60f8203c", -- 41f4
		x"000000f8", -- 41f8
		x"9c8026d8", -- 41fc
		x"59406efa", -- 4200
		x"48e7fff8", -- 4204
		x"2f052f06", -- 4208
		x"2f0b4227", -- 420c
		x"61002ce4", -- 4210
		x"61000f56", -- 4214
		x"61002cf0", -- 4218
		x"4cdf1fff", -- 421c
		x"dcbc0000", -- 4220
		x"00ff8cfc", -- 4224
		x"010048c6", -- 4228
		x"da862005", -- 422c
		x"5280e188", -- 4230
		x"b0adffee", -- 4234
		x"6f00ff58", -- 4238
		x"48e7fff8", -- 423c
		x"61002cb4", -- 4240
		x"61000f4e", -- 4244
		x"61002cc0", -- 4248
		x"4cdf1fff", -- 424c
		x"50c77cff", -- 4250
		x"0cade0ff", -- 4254
		x"ffff0028", -- 4258
		x"670a21ed", -- 425c
		x"0028fedc", -- 4260
		x"6000008e", -- 4264
		x"0cb8e0ff", -- 4268
		x"fffffedc", -- 426c
		x"66000082", -- 4270
		x"21fc0500", -- 4274
		x"0700fedc", -- 4278
		x"42072c3c", -- 427c
		x"e0ffffff", -- 4280
		x"266c001c", -- 4284
		x"4a936768", -- 4288
		x"2f0b2653", -- 428c
		x"51edffee", -- 4290
		x"48e7fff8", -- 4294
		x"558f3f3c", -- 4298
		x"000150e7", -- 429c
		x"486d0028", -- 42a0
		x"486dffee", -- 42a4
		x"51e76100", -- 42a8
		x"2c4a4eab", -- 42ac
		x"00006100", -- 42b0
		x"2c561b5f", -- 42b4
		x"ffea4cdf", -- 42b8
		x"1fff4a2d", -- 42bc
		x"ffee6728", -- 42c0
		x"0cade0ff", -- 42c4
		x"ffff0028", -- 42c8
		x"671e4a2d", -- 42cc
		x"ffea670c", -- 42d0
		x"21ed0028", -- 42d4
		x"fedc50c7", -- 42d8
		x"584f6014", -- 42dc
		x"bcbce0ff", -- 42e0
		x"ffff6604", -- 42e4
		x"2c2d0028", -- 42e8
		x"265f588b", -- 42ec
		x"d7d36094", -- 42f0
		x"206dfff2", -- 42f4
		x"21c8fdbc", -- 42f8
		x"4a07660c", -- 42fc
		x"0c86e0ff", -- 4300
		x"ffff6704", -- 4304
		x"21c6fedc", -- 4308
		x"2678fed4", -- 430c
		x"d7eb002c", -- 4310
		x"21cbfdce", -- 4314
		x"286d0024", -- 4318
		x"4240101c", -- 431c
		x"16c016dc", -- 4320
		x"53406efa", -- 4324
		x"2878fdce", -- 4328
		x"47f8fdc2", -- 432c
		x"4240101c", -- 4330
		x"32000c40", -- 4334
		x"000a6f02", -- 4338
		x"700a16dc", -- 433c
		x"53406efa", -- 4340
		x"b27c000a", -- 4344
		x"6c7416fc", -- 4348
		x"00205241", -- 434c
		x"60f26100", -- 4350
		x"2bb6588f", -- 4354
		x"21dffffc", -- 4358
		x"4e5d4cdf", -- 435c
		x"19e12f57", -- 4360
		x"0008508f", -- 4364
		x"4e756100", -- 4368
		x"2b9e0c6d", -- 436c
		x"0007fffe", -- 4370
		x"672e302d", -- 4374
		x"fffe2078", -- 4378
		x"fed42228", -- 437c
		x"005e41f8", -- 4380
		x"fdd210fc", -- 4384
		x"00206100", -- 4388
		x"1eee6100", -- 438c
		x"1f944218", -- 4390
		x"41f8fdd2", -- 4394
		x"70136018", -- 4398
		x"41fa1711", -- 439c
		x"7014600a", -- 43a0
		x"61002b64", -- 43a4
		x"41fa16f2", -- 43a8
		x"701521ed", -- 43ac
		x"ffe4fffc", -- 43b0
		x"61000a7e", -- 43b4
		x"61001412", -- 43b8
		x"60fe6100", -- 43bc
		x"caae31fc", -- 43c0
		x"4ef9ff94", -- 43c4
		x"21fc0000", -- 43c8
		x"43d2ff96", -- 43cc
		x"4e40007c", -- 43d0
		x"07002278", -- 43d4
		x"fed44ea9", -- 43d8
		x"00306100", -- 43dc
		x"30b04a29", -- 43e0
		x"00a66b18", -- 43e4
		x"286900a2", -- 43e8
		x"0c290004", -- 43ec
		x"00a66606", -- 43f0
		x"99fc0000", -- 43f4
		x"400008ac", -- 43f8
		x"00070003", -- 43fc
		x"42800838", -- 4400
		x"0003fed2", -- 4404
		x"67064aa9", -- 4408
		x"00b2671e", -- 440c
		x"246900aa", -- 4410
		x"266900ae", -- 4414
		x"725f6100", -- 4418
		x"20dc6100", -- 441c
		x"207c203c", -- 4420
		x"000000c8", -- 4424
		x"610020de", -- 4428
		x"67f443f8", -- 442c
		x"fee04280", -- 4430
		x"2878fed4", -- 4434
		x"08ac0002", -- 4438
		x"000a08ac", -- 443c
		x"0000000a", -- 4440
		x"082c0006", -- 4444
		x"000b6710", -- 4448
		x"b2fcff3a", -- 444c
		x"6706b2fc", -- 4450
		x"ffd06604", -- 4454
		x"5c89600a", -- 4458
		x"32fc4eb9", -- 445c
		x"22fc0000", -- 4460
		x"4d7ab089", -- 4464
		x"66da4ff8", -- 4468
		x"fdac1c38", -- 446c
		x"fed24e90", -- 4470
		x"600007a4", -- 4474
		x"60000010", -- 4478
		x"60000012", -- 447c
		x"60000018", -- 4480
		x"6000001c", -- 4484
		x"4e7551ef", -- 4488
		x"00044e75", -- 448c
		x"2057defc", -- 4490
		x"001451d7", -- 4494
		x"4ed02057", -- 4498
		x"defc0012", -- 449c
		x"4ed0205f", -- 44a0
		x"225f45fa", -- 44a4
		x"000e12da", -- 44a8
		x"66fc2ebc", -- 44ac
		x"000008d8", -- 44b0
		x"4ed00755", -- 44b4
		x"4e4b4e4f", -- 44b8
		x"574e0000", -- 44bc
		x"205f225f", -- 44c0
		x"12da66fc", -- 44c4
		x"4ed045fa", -- 44c8
		x"000460f0", -- 44cc
		x"05455052", -- 44d0
		x"4f4d0000", -- 44d4
		x"225f221f", -- 44d8
		x"241f205f", -- 44dc
		x"2f092278", -- 44e0
		x"fed42269", -- 44e4
		x"009ad2fc", -- 44e8
		x"00122601", -- 44ec
		x"86fc0040", -- 44f0
		x"48c3e38b", -- 44f4
		x"d3c3e189", -- 44f8
		x"d3c12009", -- 44fc
		x"0280ffff", -- 4500
		x"c000d0bc", -- 4504
		x"00004000", -- 4508
		x"9089b480", -- 450c
		x"62022002", -- 4510
		x"48e7a0c0", -- 4514
		x"4eb8315a", -- 4518
		x"4cdf0305", -- 451c
		x"94806308", -- 4520
		x"d1c0d3c0", -- 4524
		x"544960d2", -- 4528
		x"4e752078", -- 452c
		x"fed41028", -- 4530
		x"005f72ff", -- 4534
		x"2f38fffc", -- 4538
		x"3f38fffa", -- 453c
		x"31fc4ef9", -- 4540
		x"fffa21fc", -- 4544
		x"00004574", -- 4548
		x"fffc244f", -- 454c
		x"217c0002", -- 4550
		x"0000009a", -- 4554
		x"2268009a", -- 4558
		x"b3fc0040", -- 455c
		x"0000642c", -- 4560
		x"0c51f0ff", -- 4564
		x"670e06a8", -- 4568
		x"00004000", -- 456c
		x"009a60e4", -- 4570
		x"2e4a60f2", -- 4574
		x"08290003", -- 4578
		x"000367ea", -- 457c
		x"5241b001", -- 4580
		x"66e431df", -- 4584
		x"fffa21df", -- 4588
		x"fffc4e75", -- 458c
		x"31dffffa", -- 4590
		x"21dffffc", -- 4594
		x"3b7c0001", -- 4598
		x"fffe2e6d", -- 459c
		x"fff64e75", -- 45a0
		x"60004450", -- 45a4
		x"600045b2", -- 45a8
		x"60004488", -- 45ac
		x"600045aa", -- 45b0
		x"60000018", -- 45b4
		x"60000026", -- 45b8
		x"6000fedc", -- 45bc
		x"600000e8", -- 45c0
		x"4e756000", -- 45c4
		x"00fc6000", -- 45c8
		x"013c2878", -- 45cc
		x"fed4297c", -- 45d0
		x"00020000", -- 45d4
		x"006250ef", -- 45d8
		x"00044e75", -- 45dc
		x"2f38fffc", -- 45e0
		x"21fc0000", -- 45e4
		x"4694fffc", -- 45e8
		x"244f2878", -- 45ec
		x"fed4206c", -- 45f0
		x"0062b1fc", -- 45f4
		x"00400000", -- 45f8
		x"6400009c", -- 45fc
		x"0c50f0ff", -- 4600
		x"660e0c68", -- 4604
		x"f0ff0002", -- 4608
		x"67060c50", -- 460c
		x"f0ff670a", -- 4610
		x"06ac0000", -- 4614
		x"40000062", -- 4618
		x"60d40828", -- 461c
		x"00000003", -- 4620
		x"67ee1028", -- 4624
		x"000e0838", -- 4628
		x"0000fed2", -- 462c
		x"67080800", -- 4630
		x"000667dc", -- 4634
		x"60080800", -- 4638
		x"00036602", -- 463c
		x"60d2226f", -- 4640
		x"00140c11", -- 4644
		x"00016640", -- 4648
		x"10290001", -- 464c
		x"b0280002", -- 4650
		x"66be12bc", -- 4654
		x"00021368", -- 4658
		x"00020001", -- 465c
		x"42290002", -- 4660
		x"226f000c", -- 4664
		x"4291226f", -- 4668
		x"001041e8", -- 466c
		x"0008d1d0", -- 4670
		x"228843ef", -- 4674
		x"000832bc", -- 4678
		x"e94206ac", -- 467c
		x"00004000", -- 4680
		x"006250ef", -- 4684
		x"00186012", -- 4688
		x"4a290002", -- 468c
		x"67ba60c2", -- 4690
		x"2e4a6000", -- 4694
		x"ff7c51ef", -- 4698
		x"001821df", -- 469c
		x"fffc205f", -- 46a0
		x"defc0010", -- 46a4
		x"4ed0205f", -- 46a8
		x"225f45fa", -- 46ac
		x"000e12da", -- 46b0
		x"66fc2ebc", -- 46b4
		x"000008d8", -- 46b8
		x"4ed00352", -- 46bc
		x"4f4d0000", -- 46c0
		x"206f0006", -- 46c4
		x"50d0206f", -- 46c8
		x"000a20bc", -- 46cc
		x"e0ffffff", -- 46d0
		x"2078fed4", -- 46d4
		x"217ce0ff", -- 46d8
		x"ffff005e", -- 46dc
		x"558f6100", -- 46e0
		x"feea548f", -- 46e4
		x"51ef0012", -- 46e8
		x"4a2f000e", -- 46ec
		x"670c0c6f", -- 46f0
		x"00010010", -- 46f4
		x"660450ef", -- 46f8
		x"00122f57", -- 46fc
		x"000edefc", -- 4700
		x"000e4e75", -- 4704
		x"4e55fffa", -- 4708
		x"558f2f2d", -- 470c
		x"0008486d", -- 4710
		x"fffc486d", -- 4714
		x"fffc3b7c", -- 4718
		x"e942fffa", -- 471c
		x"486dfffa", -- 4720
		x"6100feba", -- 4724
		x"1b5f000c", -- 4728
		x"4e5d2f57", -- 472c
		x"0004588f", -- 4730
		x"4e756000", -- 4734
		x"4fb46000", -- 4738
		x"517c6000", -- 473c
		x"54a66000", -- 4740
		x"00166000", -- 4744
		x"56286000", -- 4748
		x"56546000", -- 474c
		x"5c966000", -- 4750
		x"583e6000", -- 4754
		x"5c8e205f", -- 4758
		x"225f45fa", -- 475c
		x"000e12da", -- 4760
		x"66fc2ebc", -- 4764
		x"00004776", -- 4768
		x"4ed00652", -- 476c
		x"454d4f54", -- 4770
		x"45001f00", -- 4774
		x"60007192", -- 4778
		x"6000765c", -- 477c
		x"60007d5e", -- 4780
		x"60000016", -- 4784
		x"60007f24", -- 4788
		x"60003a08", -- 478c
		x"60003a08", -- 4790
		x"60003a08", -- 4794
		x"60003a00", -- 4798
		x"205f225f", -- 479c
		x"45fa000e", -- 47a0
		x"12da66fc", -- 47a4
		x"2ebc0000", -- 47a8
		x"47b54ed0", -- 47ac
		x"034c414e", -- 47b0
		x"0059004d", -- 47b4
		x"41550043", -- 47b8
		x"41424c45", -- 47bc
		x"004e4f20", -- 47c0
		x"48454152", -- 47c4
		x"54424541", -- 47c8
		x"540048e7", -- 47cc
		x"64244e55", -- 47d0
		x"fffa2f09", -- 47d4
		x"42272f0a", -- 47d8
		x"486dfffa", -- 47dc
		x"4eb90000", -- 47e0
		x"d78a4a1f", -- 47e4
		x"225f6770", -- 47e8
		x"12fc002c", -- 47ec
		x"12fc0020", -- 47f0
		x"202dfffa", -- 47f4
		x"610002c0", -- 47f8
		x"302dfffe", -- 47fc
		x"610002c6", -- 4800
		x"4e5d42a7", -- 4804
		x"2f0a42a7", -- 4808
		x"4eb90000", -- 480c
		x"d7cc4a9f", -- 4810
		x"66722a78", -- 4814
		x"fed4082d", -- 4818
		x"0000000a", -- 481c
		x"673e42a7", -- 4820
		x"2f0a2f3c", -- 4824
		x"00000001", -- 4828
		x"4eb90000", -- 482c
		x"d7cc241f", -- 4830
		x"672a45fa", -- 4834
		x"ff7f0c02", -- 4838
		x"001b6724", -- 483c
		x"45faff79", -- 4840
		x"0c020019", -- 4844
		x"671a0c02", -- 4848
		x"001a6714", -- 484c
		x"45faff6f", -- 4850
		x"0c020023", -- 4854
		x"670a602c", -- 4858
		x"4e5d6028", -- 485c
		x"51c06026", -- 4860
		x"421141f8", -- 4864
		x"fdd26100", -- 4868
		x"0f1443f8", -- 486c
		x"fdd222fc", -- 4870
		x"20202020", -- 4874
		x"12da66fc", -- 4878
		x"93fc0000", -- 487c
		x"00010c02", -- 4880
		x"002367d8", -- 4884
		x"50c04cdf", -- 4888
		x"24264e75", -- 488c
		x"4238fdcd", -- 4890
		x"4e7544fc", -- 4894
		x"00004e75", -- 4898
		x"2a4f0838", -- 489c
		x"0005fed2", -- 48a0
		x"662a7024", -- 48a4
		x"6100058a", -- 48a8
		x"4dfa0016", -- 48ac
		x"41f90047", -- 48b0
		x"80006122", -- 48b4
		x"4a00670c", -- 48b8
		x"41fa12ce", -- 48bc
		x"600005c2", -- 48c0
		x"2e4d4e75", -- 48c4
		x"41fa12c2", -- 48c8
		x"600005b2", -- 48cc
		x"7c036100", -- 48d0
		x"07d267ec", -- 48d4
		x"4e7543e8", -- 48d8
		x"00176100", -- 48dc
		x"009c0828", -- 48e0
		x"00070005", -- 48e4
		x"660c0828", -- 48e8
		x"00060005", -- 48ec
		x"67000082", -- 48f0
		x"60760828", -- 48f4
		x"00060005", -- 48f8
		x"66761028", -- 48fc
		x"0017c03c", -- 4900
		x"00cb5300", -- 4904
		x"666a1028", -- 4908
		x"0015c03c", -- 490c
		x"00e66660", -- 4910
		x"12bc008a", -- 4914
		x"10280015", -- 4918
		x"c03c00e6", -- 491c
		x"903c0002", -- 4920
		x"664e12bc", -- 4924
		x"00891028", -- 4928
		x"0015c03c", -- 492c
		x"00e6b03c", -- 4930
		x"0084663c", -- 4934
		x"12bc0009", -- 4938
		x"12bc000c", -- 493c
		x"727f4a28", -- 4940
		x"00175bc9", -- 4944
		x"fffa6a28", -- 4948
		x"10280015", -- 494c
		x"c03c00e6", -- 4950
		x"b03c00a0", -- 4954
		x"661a0108", -- 4958
		x"00110240", -- 495c
		x"fffdb07c", -- 4960
		x"1200660c", -- 4964
		x"12bc000b", -- 4968
		x"51c012bc", -- 496c
		x"00104e75", -- 4970
		x"50c012bc", -- 4974
		x"00104e75", -- 4978
		x"12bc0080", -- 497c
		x"12bc0093", -- 4980
		x"70000188", -- 4984
		x"00111028", -- 4988
		x"0005b1fc", -- 498c
		x"00478000", -- 4990
		x"660c0800", -- 4994
		x"00076704", -- 4998
		x"70156002", -- 499c
		x"70140240", -- 49a0
		x"001f0c40", -- 49a4
		x"001f6602", -- 49a8
		x"70001140", -- 49ac
		x"001912bc", -- 49b0
		x"00000828", -- 49b4
		x"00070005", -- 49b8
		x"671c12bc", -- 49bc
		x"001012bc", -- 49c0
		x"008f4878", -- 49c4
		x"00646100", -- 49c8
		x"60c212bc", -- 49cc
		x"000f12bc", -- 49d0
		x"009012bc", -- 49d4
		x"000b4e75", -- 49d8
		x"4dfa003e", -- 49dc
		x"117c0080", -- 49e0
		x"0016117c", -- 49e4
		x"00000012", -- 49e8
		x"117c0007", -- 49ec
		x"0010117c", -- 49f0
		x"00070016", -- 49f4
		x"117c001f", -- 49f8
		x"00181a3c", -- 49fc
		x"00011145", -- 4a00
		x"00104878", -- 4a04
		x"03e86100", -- 4a08
		x"6082ba28", -- 4a0c
		x"00106608", -- 4a10
		x"e30d64ea", -- 4a14
		x"51c06002", -- 4a18
		x"50c04dfa", -- 4a1c
		x"001a117c", -- 4a20
		x"00000018", -- 4a24
		x"117c0080", -- 4a28
		x"0016117c", -- 4a2c
		x"00400010", -- 4a30
		x"117c0007", -- 4a34
		x"00164e75", -- 4a38
		x"4dfa0022", -- 4a3c
		x"2a4f117c", -- 4a40
		x"00000001", -- 4a44
		x"61002df0", -- 4a48
		x"2a48dbfc", -- 4a4c
		x"00008000", -- 4a50
		x"2248d3fc", -- 4a54
		x"00020000", -- 4a58
		x"60000530", -- 4a5c
		x"2e4d50c0", -- 4a60
		x"4e756100", -- 4a64
		x"373a0838", -- 4a68
		x"0006feda", -- 4a6c
		x"661641fa", -- 4a70
		x"121d0838", -- 4a74
		x"0000fed9", -- 4a78
		x"66066100", -- 4a7c
		x"04006004", -- 4a80
		x"610003fe", -- 4a84
		x"4e75780a", -- 4a88
		x"22006a06", -- 4a8c
		x"12fc002d", -- 4a90
		x"44813401", -- 4a94
		x"42414841", -- 4a98
		x"82c43601", -- 4a9c
		x"320282c4", -- 4aa0
		x"34013203", -- 4aa4
		x"48413f01", -- 4aa8
		x"86426702", -- 4aac
		x"61e67230", -- 4ab0
		x"d25f12c1", -- 4ab4
		x"4e754840", -- 4ab8
		x"610a4840", -- 4abc
		x"60064840", -- 4ac0
		x"610a4840", -- 4ac4
		x"3200e058", -- 4ac8
		x"61023001", -- 4acc
		x"3400e850", -- 4ad0
		x"61023002", -- 4ad4
		x"0200000f", -- 4ad8
		x"00000030", -- 4adc
		x"0c000039", -- 4ae0
		x"6f025e40", -- 4ae4
		x"12c04e75", -- 4ae8
		x"12d866fc", -- 4aec
		x"53894e75", -- 4af0
		x"48e780c0", -- 4af4
		x"31fc4ef9", -- 4af8
		x"ff5821fc", -- 4afc
		x"00004c14", -- 4b00
		x"ff5a41f8", -- 4b04
		x"ff5e43f8", -- 4b08
		x"ff9a30fc", -- 4b0c
		x"4ef920fc", -- 4b10
		x"00004c0e", -- 4b14
		x"b3c862f2", -- 4b18
		x"5c4843f8", -- 4b1c
		x"ffbe0c50", -- 4b20
		x"4ef96604", -- 4b24
		x"5c48600a", -- 4b28
		x"30fc4eb9", -- 4b2c
		x"20fc0000", -- 4b30
		x"4db8b3c8", -- 4b34
		x"62e84280", -- 4b38
		x"43f8ffd0", -- 4b3c
		x"41f8ffc4", -- 4b40
		x"30fc4ef9", -- 4b44
		x"20fc0000", -- 4b48
		x"4c0eb3c8", -- 4b4c
		x"62f25c48", -- 4b50
		x"30fc4ef9", -- 4b54
		x"20fc0000", -- 4b58
		x"4c0eb1c0", -- 4b5c
		x"66e24cdf", -- 4b60
		x"03014e75", -- 4b64
		x"2878fed4", -- 4b68
		x"206c0010", -- 4b6c
		x"30f8ff58", -- 4b70
		x"20f8ff5a", -- 4b74
		x"49f8ff76", -- 4b78
		x"20dc20dc", -- 4b7c
		x"20dc31fc", -- 4b80
		x"4ef9ff58", -- 4b84
		x"21fc0000", -- 4b88
		x"4c14ff5a", -- 4b8c
		x"31fc4ef9", -- 4b90
		x"ff7c21fc", -- 4b94
		x"00004c0e", -- 4b98
		x"ff7e31fc", -- 4b9c
		x"4ef9ff76", -- 4ba0
		x"21fc0000", -- 4ba4
		x"4c0eff78", -- 4ba8
		x"4e752878", -- 4bac
		x"fed4206c", -- 4bb0
		x"001031d8", -- 4bb4
		x"ff5821d8", -- 4bb8
		x"ff5a49f8", -- 4bbc
		x"ff7628d8", -- 4bc0
		x"28d828d8", -- 4bc4
		x"4e75bffc", -- 4bc8
		x"00000100", -- 4bcc
		x"63044ef8", -- 4bd0
		x"fffa4ff8", -- 4bd4
		x"01004ed6", -- 4bd8
		x"4ebac3ee", -- 4bdc
		x"4ed64e73", -- 4be0
		x"31fc4ef9", -- 4be4
		x"fffa21fc", -- 4be8
		x"00004bdc", -- 4bec
		x"fffc4e75", -- 4bf0
		x"31fc4ef9", -- 4bf4
		x"ff9a21fc", -- 4bf8
		x"00004be2", -- 4bfc
		x"ff9c6004", -- 4c00
		x"4e722600", -- 4c04
		x"4e722700", -- 4c08
		x"60fa3b7c", -- 4c0c
		x"0006fffe", -- 4c10
		x"2e6dfff6", -- 4c14
		x"4e753f38", -- 4c18
		x"fffa2f38", -- 4c1c
		x"fffc31fc", -- 4c20
		x"4ef9fffa", -- 4c24
		x"21fc0000", -- 4c28
		x"4c4efffc", -- 4c2c
		x"6100c274", -- 4c30
		x"0c794ef9", -- 4c34
		x"00880000", -- 4c38
		x"661421df", -- 4c3c
		x"fffc31df", -- 4c40
		x"fffa6100", -- 4c44
		x"c25e588f", -- 4c48
		x"4e754eba", -- 4c4c
		x"c37c21df", -- 4c50
		x"fffc31df", -- 4c54
		x"fffa6100", -- 4c58
		x"c24a4e75", -- 4c5c
		x"48e7fffe", -- 4c60
		x"4dfa0064", -- 4c64
		x"3039005b", -- 4c68
		x"00004279", -- 4c6c
		x"005b0000", -- 4c70
		x"b1f8fdd2", -- 4c74
		x"660a33fc", -- 4c78
		x"0001005b", -- 4c7c
		x"00006046", -- 4c80
		x"6100c1e8", -- 4c84
		x"200821c8", -- 4c88
		x"fdd2b290", -- 4c8c
		x"670641fa", -- 4c90
		x"0f8f6004", -- 4c94
		x"41fa0f9f", -- 4c98
		x"43f8fdd6", -- 4c9c
		x"6100fe4a", -- 4ca0
		x"6100fe14", -- 4ca4
		x"421941f8", -- 4ca8
		x"fdd66100", -- 4cac
		x"0ad021fc", -- 4cb0
		x"00004cde", -- 4cb4
		x"ff244cdf", -- 4cb8
		x"7fff33fc", -- 4cbc
		x"0001005b", -- 4cc0
		x"0000b290", -- 4cc4
		x"60064cdf", -- 4cc8
		x"7fff4e73", -- 4ccc
		x"21fc0000", -- 4cd0
		x"4c60ff24", -- 4cd4
		x"6100c1b6", -- 4cd8
		x"4e7348e7", -- 4cdc
		x"fffe4dfa", -- 4ce0
		x"ffe63039", -- 4ce4
		x"005b0000", -- 4ce8
		x"4279005b", -- 4cec
		x"00002878", -- 4cf0
		x"fed411ec", -- 4cf4
		x"000afdd6", -- 4cf8
		x"4cdf7fff", -- 4cfc
		x"76007801", -- 4d00
		x"08380000", -- 4d04
		x"fdd66706", -- 4d08
		x"4be80004", -- 4d0c
		x"600449e8", -- 4d10
		x"000433fc", -- 4d14
		x"0001005b", -- 4d18
		x"00004e73", -- 4d1c
		x"bffc0000", -- 4d20
		x"0100634e", -- 4d24
		x"08380003", -- 4d28
		x"fed26628", -- 4d2c
		x"08390002", -- 4d30
		x"00478005", -- 4d34
		x"673c48e7", -- 4d38
		x"00602278", -- 4d3c
		x"fed42469", -- 4d40
		x"00aa0812", -- 4d44
		x"00024cdf", -- 4d48
		x"06006604", -- 4d4c
		x"4ef8ff34", -- 4d50
		x"4ef8ff2e", -- 4d54
		x"48e70060", -- 4d58
		x"2278fed4", -- 4d5c
		x"4aa900b2", -- 4d60
		x"67102469", -- 4d64
		x"00b2082a", -- 4d68
		x"00030003", -- 4d6c
		x"66d04cdf", -- 4d70
		x"06004ef8", -- 4d74
		x"ff2221d7", -- 4d78
		x"fdbc31fc", -- 4d7c
		x"4ef9ff94", -- 4d80
		x"21fc0000", -- 4d84
		x"4d8eff96", -- 4d88
		x"4e402078", -- 4d8c
		x"fed44ea8", -- 4d90
		x"003043f8", -- 4d94
		x"fdd241fa", -- 4d98
		x"0cec6100", -- 4d9c
		x"fd4c2038", -- 4da0
		x"fdbc5d80", -- 4da4
		x"6100fd10", -- 4da8
		x"421941f8", -- 4dac
		x"fdd26100", -- 4db0
		x"0a1860fe", -- 4db4
		x"21d7fdbc", -- 4db8
		x"60d82f0e", -- 4dbc
		x"4dfa0008", -- 4dc0
		x"10390044", -- 4dc4
		x"c00031fc", -- 4dc8
		x"4eb9ffb8", -- 4dcc
		x"21fc0000", -- 4dd0
		x"4db8ffba", -- 4dd4
		x"2c5f4e73", -- 4dd8
		x"08f80000", -- 4ddc
		x"fdcc4e75", -- 4de0
		x"3b7c0820", -- 4de4
		x"fffe6000", -- 4de8
		x"00083b7c", -- 4dec
		x"0820fffe", -- 4df0
		x"2e6dfff6", -- 4df4
		x"4e753b7c", -- 4df8
		x"0820fffe", -- 4dfc
		x"60f23b7c", -- 4e00
		x"0820fffe", -- 4e04
		x"60ea2078", -- 4e08
		x"fed4217c", -- 4e0c
		x"fffffac0", -- 4e10
		x"03302238", -- 4e14
		x"fed47020", -- 4e18
		x"c0e80334", -- 4e1c
		x"d28021c1", -- 4e20
		x"fdce2028", -- 4e24
		x"0014d1b8", -- 4e28
		x"fdce2141", -- 4e2c
		x"00104e75", -- 4e30
		x"48e78008", -- 4e34
		x"2878fed4", -- 4e38
		x"1940009e", -- 4e3c
		x"4a6c00a0", -- 4e40
		x"6b084600", -- 4e44
		x"13c00001", -- 4e48
		x"ffff4cdf", -- 4e4c
		x"10014e75", -- 4e50
		x"48e7e008", -- 4e54
		x"2878fed4", -- 4e58
		x"102c009e", -- 4e5c
		x"122c00a1", -- 4e60
		x"67100c00", -- 4e64
		x"0010670a", -- 4e68
		x"0c010010", -- 4e6c
		x"6708b001", -- 4e70
		x"62041940", -- 4e74
		x"00a14cdf", -- 4e78
		x"10074e75", -- 4e7c
		x"600008fe", -- 4e80
		x"48e700c0", -- 4e84
		x"61ca43f8", -- 4e88
		x"fdd212d8", -- 4e8c
		x"66fc5349", -- 4e90
		x"41fa0dc6", -- 4e94
		x"12d866fc", -- 4e98
		x"41f8fdd2", -- 4e9c
		x"610008de", -- 4ea0
		x"4cdf0300", -- 4ea4
		x"4e757200", -- 4ea8
		x"74007600", -- 4eac
		x"0b080000", -- 4eb0
		x"0d080001", -- 4eb4
		x"d445d541", -- 4eb8
		x"d646d741", -- 4ebc
		x"58485984", -- 4ec0
		x"6eea5242", -- 4ec4
		x"30025243", -- 4ec8
		x"8043bffc", -- 4ecc
		x"00000100", -- 4ed0
		x"63024e75", -- 4ed4
		x"4ed47200", -- 4ed8
		x"74007600", -- 4edc
		x"0b080000", -- 4ee0
		x"0d080001", -- 4ee4
		x"4206d445", -- 4ee8
		x"d541d646", -- 4eec
		x"d7415848", -- 4ef0
		x"59846eb8", -- 4ef4
		x"60d4e318", -- 4ef8
		x"e158e318", -- 4efc
		x"e1584840", -- 4f00
		x"4e75204a", -- 4f04
		x"223cee11", -- 4f08
		x"ee1103c8", -- 4f0c
		x"00005088", -- 4f10
		x"b3c866f6", -- 4f14
		x"76ff78ff", -- 4f18
		x"4dfa0060", -- 4f1c
		x"74fe203c", -- 4f20
		x"ee11ee11", -- 4f24
		x"223c8877", -- 4f28
		x"88775242", -- 4f2c
		x"c14161c6", -- 4f30
		x"61c42a01", -- 4f34
		x"ca870802", -- 4f38
		x"0001661e", -- 4f3c
		x"20495188", -- 4f40
		x"0d480000", -- 4f44
		x"cc87ba86", -- 4f48
		x"662801c8", -- 4f4c
		x"0000b1ca", -- 4f50
		x"62ec0c00", -- 4f54
		x"001166d2", -- 4f58
		x"602c204a", -- 4f5c
		x"0d480000", -- 4f60
		x"cc87ba86", -- 4f64
		x"660c01c8", -- 4f68
		x"00005088", -- 4f6c
		x"b1c966ec", -- 4f70
		x"60e02605", -- 4f74
		x"09480000", -- 4f78
		x"c8872478", -- 4f7c
		x"fed42548", -- 4f80
		x"032870ff", -- 4f84
		x"4e754240", -- 4f88
		x"4e754dfa", -- 4f8c
		x"0038203c", -- 4f90
		x"eeee1111", -- 4f94
		x"22002401", -- 4f98
		x"26022803", -- 4f9c
		x"2a042c05", -- 4fa0
		x"2e062049", -- 4fa4
		x"48e0ff00", -- 4fa8
		x"b1cd62f8", -- 4fac
		x"76ff78ff", -- 4fb0
		x"264d6100", -- 4fb4
		x"b6a8bbcb", -- 4fb8
		x"670e598d", -- 4fbc
		x"2078fed4", -- 4fc0
		x"214d0328", -- 4fc4
		x"50c04e75", -- 4fc8
		x"51c04e75", -- 4fcc
		x"48e7fffe", -- 4fd0
		x"2878fed4", -- 4fd4
		x"08380003", -- 4fd8
		x"fed26706", -- 4fdc
		x"4aac00b2", -- 4fe0
		x"67327606", -- 4fe4
		x"38002878", -- 4fe8
		x"fed4082c", -- 4fec
		x"0002005c", -- 4ff0
		x"67220704", -- 4ff4
		x"6706343c", -- 4ff8
		x"10cd6004", -- 4ffc
		x"343c04cd", -- 5000
		x"61001886", -- 5004
		x"4dfab8ce", -- 5008
		x"303c03e8", -- 500c
		x"61002c04", -- 5010
		x"53436cd2", -- 5014
		x"4cdf7fff", -- 5018
		x"4e75b883", -- 501c
		x"676848e7", -- 5020
		x"fffe43f8", -- 5024
		x"fdd241fa", -- 5028
		x"0bd54a83", -- 502c
		x"6708b883", -- 5030
		x"660441fa", -- 5034
		x"0bdb6100", -- 5038
		x"fab02078", -- 503c
		x"fed42028", -- 5040
		x"03286100", -- 5044
		x"fa724219", -- 5048
		x"41f8fdd2", -- 504c
		x"6100072e", -- 5050
		x"4a83672e", -- 5054
		x"b883672a", -- 5058
		x"43f8fdd2", -- 505c
		x"22fc2028", -- 5060
		x"573a2003", -- 5064
		x"6100fa50", -- 5068
		x"22fc2c20", -- 506c
		x"523a2004", -- 5070
		x"6100fa44", -- 5074
		x"12fc0029", -- 5078
		x"421941f8", -- 507c
		x"fdd26100", -- 5080
		x"06fc4cdf", -- 5084
		x"7fff4e75", -- 5088
		x"41fa0a4f", -- 508c
		x"611041fa", -- 5090
		x"0a59610a", -- 5094
		x"41fa0a6c", -- 5098
		x"610441fa", -- 509c
		x"0a7b6000", -- 50a0
		x"06dc70ff", -- 50a4
		x"4e75203c", -- 50a8
		x"ffffc000", -- 50ac
		x"b9c06304", -- 50b0
		x"70ff4e75", -- 50b4
		x"70004e75", -- 50b8
		x"48a7c000", -- 50bc
		x"2078fed4", -- 50c0
		x"1028005e", -- 50c4
		x"12000201", -- 50c8
		x"00e00c01", -- 50cc
		x"00e06702", -- 50d0
		x"10012068", -- 50d4
		x"00204a90", -- 50d8
		x"670ab028", -- 50dc
		x"00086704", -- 50e0
		x"d1d060f2", -- 50e4
		x"20680004", -- 50e8
		x"4c9f0003", -- 50ec
		x"4e754ef9", -- 50f0
		x"000101d6", -- 50f4
		x"4ef90001", -- 50f8
		x"000e2078", -- 50fc
		x"fed4216f", -- 5100
		x"0004005e", -- 5104
		x"2f570004", -- 5108
		x"588f6100", -- 510c
		x"fa584e55", -- 5110
		x"fff6487a", -- 5114
		x"001a2b4f", -- 5118
		x"fff6554f", -- 511c
		x"619a4ea8", -- 5120
		x"00003b57", -- 5124
		x"00086100", -- 5128
		x"fa824e5d", -- 512c
		x"4e756100", -- 5130
		x"fa7a302d", -- 5134
		x"fffe4e5d", -- 5138
		x"3b40fffe", -- 513c
		x"2e6dfff6", -- 5140
		x"4e756100", -- 5144
		x"fa204cdf", -- 5148
		x"001f2f00", -- 514c
		x"4e55fff6", -- 5150
		x"487affdc", -- 5154
		x"2b4ffff6", -- 5158
		x"554f48e7", -- 515c
		x"78006100", -- 5160
		x"ff584ea8", -- 5164
		x"000460ba", -- 5168
		x"6100f9fa", -- 516c
		x"4cdf000f", -- 5170
		x"381f2f00", -- 5174
		x"4e55fff6", -- 5178
		x"487affb4", -- 517c
		x"2b4ffff6", -- 5180
		x"3f0448e7", -- 5184
		x"70006100", -- 5188
		x"ff304ea8", -- 518c
		x"00086096", -- 5190
		x"6100f9d2", -- 5194
		x"4e55fff6", -- 5198
		x"487aff94", -- 519c
		x"2b4ffff6", -- 51a0
		x"6100ff16", -- 51a4
		x"4ea80010", -- 51a8
		x"6000ff7c", -- 51ac
		x"6100ff0a", -- 51b0
		x"4ee8000c", -- 51b4
		x"600035c6", -- 51b8
		x"6000399e", -- 51bc
		x"600036d0", -- 51c0
		x"60003996", -- 51c4
		x"600038e8", -- 51c8
		x"6000398e", -- 51cc
		x"60003922", -- 51d0
		x"60003986", -- 51d4
		x"41f9005f", -- 51d8
		x"80000148", -- 51dc
		x"00090348", -- 51e0
		x"0009b181", -- 51e4
		x"48414a41", -- 51e8
		x"67044841", -- 51ec
		x"b3804e75", -- 51f0
		x"48e78080", -- 51f4
		x"206f000c", -- 51f8
		x"2f6f0008", -- 51fc
		x"000c2010", -- 5200
		x"ed889090", -- 5204
		x"e3889090", -- 5208
		x"e78890bc", -- 520c
		x"00000019", -- 5210
		x"20804cdf", -- 5214
		x"0101588f", -- 5218
		x"4e7548e7", -- 521c
		x"c08061b4", -- 5220
		x"206f0010", -- 5224
		x"221092bc", -- 5228
		x"00000010", -- 522c
		x"e4899081", -- 5230
		x"20804cdf", -- 5234
		x"01032e9f", -- 5238
		x"4e7548e7", -- 523c
		x"c0806194", -- 5240
		x"206f0010", -- 5244
		x"2f6f000c", -- 5248
		x"0010b090", -- 524c
		x"4cdf0103", -- 5250
		x"588f4e75", -- 5254
		x"422f0008", -- 5258
		x"2f2f0004", -- 525c
		x"61dc6a06", -- 5260
		x"1f7c0001", -- 5264
		x"00082e9f", -- 5268
		x"4e7548e7", -- 526c
		x"c08041f9", -- 5270
		x"005f8000", -- 5274
		x"01480009", -- 5278
		x"03480009", -- 527c
		x"b1814841", -- 5280
		x"4a416704", -- 5284
		x"4841b380", -- 5288
		x"222f0010", -- 528c
		x"e4895b81", -- 5290
		x"6f0a9081", -- 5294
		x"03480009", -- 5298
		x"b2806af8", -- 529c
		x"4cdf0103", -- 52a0
		x"2e9f4e75", -- 52a4
		x"48e7fcf8", -- 52a8
		x"2078fed4", -- 52ac
		x"1a28000b", -- 52b0
		x"74046106", -- 52b4
		x"4cdf1f3f", -- 52b8
		x"4e752078", -- 52bc
		x"fed44aa8", -- 52c0
		x"00486708", -- 52c4
		x"610000d4", -- 52c8
		x"600000c4", -- 52cc
		x"08380004", -- 52d0
		x"fed26716", -- 52d4
		x"30390051", -- 52d8
		x"fffe0800", -- 52dc
		x"000f6600", -- 52e0
		x"00a4e648", -- 52e4
		x"c07c001f", -- 52e8
		x"602e0838", -- 52ec
		x"0005fed2", -- 52f0
		x"660e0839", -- 52f4
		x"00020047", -- 52f8
		x"80036704", -- 52fc
		x"70046018", -- 5300
		x"42400805", -- 5304
		x"00076620", -- 5308
		x"08380000", -- 530c
		x"fed26618", -- 5310
		x"70023239", -- 5314
		x"00512704", -- 5318
		x"08800000", -- 531c
		x"08050000", -- 5320
		x"671008c0", -- 5324
		x"0000600a", -- 5328
		x"08380000", -- 532c
		x"fed26602", -- 5330
		x"70ff41fa", -- 5334
		x"024a0c40", -- 5338
		x"000b6e52", -- 533c
		x"3200e349", -- 5340
		x"32301000", -- 5344
		x"67480805", -- 5348
		x"00076714", -- 534c
		x"08000000", -- 5350
		x"67084a39", -- 5354
		x"00514001", -- 5358
		x"60064a39", -- 535c
		x"00515001", -- 5360
		x"08000000", -- 5364
		x"67084a79", -- 5368
		x"00516000", -- 536c
		x"60064a79", -- 5370
		x"00516004", -- 5374
		x"41f01000", -- 5378
		x"720fd0c2", -- 537c
		x"924243f9", -- 5380
		x"00510001", -- 5384
		x"12811358", -- 5388
		x"000251c9", -- 538c
		x"fff8bffc", -- 5390
		x"00000100", -- 5394
		x"63024e75", -- 5398
		x"4ed42078", -- 539c
		x"fed42068", -- 53a0
		x"00484200", -- 53a4
		x"42814282", -- 53a8
		x"02280060", -- 53ac
		x"0001660c", -- 53b0
		x"12284001", -- 53b4
		x"c23c0030", -- 53b8
		x"e8497001", -- 53bc
		x"4a01660a", -- 53c0
		x"05080023", -- 53c4
		x"43f02800", -- 53c8
		x"60280c01", -- 53cc
		x"0001660a", -- 53d0
		x"05080027", -- 53d4
		x"43f02800", -- 53d8
		x"60180c01", -- 53dc
		x"0002660a", -- 53e0
		x"0508002b", -- 53e4
		x"43f02800", -- 53e8
		x"60080508", -- 53ec
		x"002f43f0", -- 53f0
		x"28004241", -- 53f4
		x"18290000", -- 53f8
		x"12290002", -- 53fc
		x"05090004", -- 5400
		x"508945f0", -- 5404
		x"28000804", -- 5408
		x"00006628", -- 540c
		x"08040006", -- 5410
		x"660e0509", -- 5414
		x"00005849", -- 5418
		x"34c251c9", -- 541c
		x"fff66054", -- 5420
		x"05090000", -- 5424
		x"07090004", -- 5428
		x"508934c2", -- 542c
		x"34c35541", -- 5430
		x"6b4260f6", -- 5434
		x"2f3c002d", -- 5438
		x"c6c04857", -- 543c
		x"6100fddc", -- 5440
		x"14290002", -- 5444
		x"02820000", -- 5448
		x"000f4a29", -- 544c
		x"00006612", -- 5450
		x"48576100", -- 5454
		x"fde66b08", -- 5458
		x"36120503", -- 545c
		x"66f26010", -- 5460
		x"4ed64857", -- 5464
		x"6100fdd4", -- 5468
		x"6bf63612", -- 546c
		x"050367f2", -- 5470
		x"584f5849", -- 5474
		x"08040007", -- 5478
		x"6700ff78", -- 547c
		x"4a00665e", -- 5480
		x"52400308", -- 5484
		x"00334a41", -- 5488
		x"67544281", -- 548c
		x"03080057", -- 5490
		x"4a41670e", -- 5494
		x"43f01800", -- 5498
		x"14110282", -- 549c
		x"00000003", -- 54a0
		x"660c0508", -- 54a4
		x"003f43f0", -- 54a8
		x"28006000", -- 54ac
		x"ff460c02", -- 54b0
		x"0001660c", -- 54b4
		x"05080043", -- 54b8
		x"43f02800", -- 54bc
		x"6000ff34", -- 54c0
		x"0c010002", -- 54c4
		x"660c0508", -- 54c8
		x"004743f0", -- 54cc
		x"28006000", -- 54d0
		x"ff220508", -- 54d4
		x"004b43f0", -- 54d8
		x"28006000", -- 54dc
		x"ff16bffc", -- 54e0
		x"00000100", -- 54e4
		x"63024e75", -- 54e8
		x"4ed448e7", -- 54ec
		x"fcf82078", -- 54f0
		x"fed44aa8", -- 54f4
		x"00486706", -- 54f8
		x"61000194", -- 54fc
		x"60780c28", -- 5500
		x"008000a6", -- 5504
		x"665a6100", -- 5508
		x"22c4606a", -- 550c
		x"48e7fcf8", -- 5510
		x"2078fed4", -- 5514
		x"1038fed2", -- 5518
		x"4aa80048", -- 551c
		x"670a6100", -- 5520
		x"fe7a6100", -- 5524
		x"017c604e", -- 5528
		x"0c280080", -- 552c
		x"00a6660a", -- 5530
		x"610022ce", -- 5534
		x"61002296", -- 5538
		x"603cc07c", -- 553c
		x"00070c40", -- 5540
		x"0002660e", -- 5544
		x"4a790051", -- 5548
		x"600433fc", -- 554c
		x"00000051", -- 5550
		x"21a02078", -- 5554
		x"fed41a28", -- 5558
		x"000b4242", -- 555c
		x"6100fd5c", -- 5560
		x"203c0020", -- 5564
		x"002041f9", -- 5568
		x"0051a000", -- 556c
		x"20c0b1fc", -- 5570
		x"0051b000", -- 5574
		x"6df64cdf", -- 5578
		x"1f3f4e75", -- 557c
		x"00280018", -- 5580
		x"00000038", -- 5584
		x"00480058", -- 5588
		x"00680078", -- 558c
		x"00880098", -- 5590
		x"00a80000", -- 5594
		x"00b88233", -- 5598
		x"82330b4b", -- 559c
		x"0b001919", -- 55a0
		x"09190a31", -- 55a4
		x"3240d030", -- 55a8
		x"d0300b4a", -- 55ac
		x"0b001919", -- 55b0
		x"0919024f", -- 55b4
		x"5067d030", -- 55b8
		x"d0300d4c", -- 55bc
		x"0e001919", -- 55c0
		x"0a1a064c", -- 55c4
		x"5072d030", -- 55c8
		x"d0300d4c", -- 55cc
		x"0e001c19", -- 55d0
		x"0320064c", -- 55d4
		x"5072d030", -- 55d8
		x"d0300b4b", -- 55dc
		x"0b001919", -- 55e0
		x"08190b4f", -- 55e4
		x"5067d030", -- 55e8
		x"d0300b4b", -- 55ec
		x"0b001e19", -- 55f0
		x"001f0b4f", -- 55f4
		x"5067d030", -- 55f8
		x"d0300d4c", -- 55fc
		x"0e001819", -- 5600
		x"0a1ae762", -- 5604
		x"5072d030", -- 5608
		x"d0300d4c", -- 560c
		x"0e001b19", -- 5610
		x"03207762", -- 5614
		x"5072d030", -- 5618
		x"d0300b4a", -- 561c
		x"0b001919", -- 5620
		x"031a0d50", -- 5624
		x"5065d030", -- 5628
		x"d0300b4a", -- 562c
		x"0b001c19", -- 5630
		x"041f1455", -- 5634
		x"5066d030", -- 5638
		x"d0300b4a", -- 563c
		x"0b001919", -- 5640
		x"03191660", -- 5644
		x"507e5240", -- 5648
		x"600000aa", -- 564c
		x"700041f9", -- 5650
		x"00538000", -- 5654
		x"323c1fff", -- 5658
		x"08380004", -- 565c
		x"fed26726", -- 5660
		x"7418c439", -- 5664
		x"0051fffe", -- 5668
		x"671c08b9", -- 566c
		x"00000051", -- 5670
		x"fffd41f9", -- 5674
		x"00520000", -- 5678
		x"72ff0839", -- 567c
		x"00030051", -- 5680
		x"fffe6602", -- 5684
		x"e24920c0", -- 5688
		x"51c9fffc", -- 568c
		x"4e7548e7", -- 5690
		x"f0c02078", -- 5694
		x"fed42068", -- 5698
		x"00480108", -- 569c
		x"00116010", -- 56a0
		x"48e7f0c0", -- 56a4
		x"2078fed4", -- 56a8
		x"20680048", -- 56ac
		x"01080009", -- 56b0
		x"240c49fa", -- 56b4
		x"00066100", -- 56b8
		x"08fa2243", -- 56bc
		x"28420508", -- 56c0
		x"0005c0c2", -- 56c4
		x"e4885380", -- 56c8
		x"243c0000", -- 56cc
		x"000022c2", -- 56d0
		x"51c8fffc", -- 56d4
		x"42405380", -- 56d8
		x"6ef4bffc", -- 56dc
		x"00000100", -- 56e0
		x"63064cdf", -- 56e4
		x"030f4e75", -- 56e8
		x"4ed448e7", -- 56ec
		x"c0c02278", -- 56f0
		x"fed46010", -- 56f4
		x"48e7c0c0", -- 56f8
		x"2278fed4", -- 56fc
		x"32007001", -- 5700
		x"4ea9003c", -- 5704
		x"42401018", -- 5708
		x"67064ea9", -- 570c
		x"003660f6", -- 5710
		x"4cdf0303", -- 5714
		x"4e7548e7", -- 5718
		x"c0082878", -- 571c
		x"fed43200", -- 5720
		x"70014eac", -- 5724
		x"003c4240", -- 5728
		x"b26c0056", -- 572c
		x"660270ff", -- 5730
		x"322c0046", -- 5734
		x"d240303c", -- 5738
		x"00204eac", -- 573c
		x"00365341", -- 5740
		x"6ef84cdf", -- 5744
		x"10034e75", -- 5748
		x"48e7e008", -- 574c
		x"2878fed4", -- 5750
		x"322c0056", -- 5754
		x"5541302c", -- 5758
		x"0046e248", -- 575c
		x"52404eac", -- 5760
		x"003c7020", -- 5764
		x"342c0046", -- 5768
		x"e24a4eac", -- 576c
		x"00365342", -- 5770
		x"6ef85341", -- 5774
		x"6ee04cdf", -- 5778
		x"10074e75", -- 577c
		x"48e7c088", -- 5780
		x"2878fed4", -- 5784
		x"7001322c", -- 5788
		x"032e4eac", -- 578c
		x"003c526c", -- 5790
		x"032e302c", -- 5794
		x"00565540", -- 5798
		x"b06c032e", -- 579c
		x"6c06397c", -- 57a0
		x"0001032e", -- 57a4
		x"322c0046", -- 57a8
		x"e2491018", -- 57ac
		x"670e4eac", -- 57b0
		x"00365341", -- 57b4
		x"6ef44cdf", -- 57b8
		x"11034e75", -- 57bc
		x"70204eac", -- 57c0
		x"00365341", -- 57c4
		x"6ef860ee", -- 57c8
		x"48e78008", -- 57cc
		x"2878fed4", -- 57d0
		x"302c0056", -- 57d4
		x"53406100", -- 57d8
		x"ff3e6100", -- 57dc
		x"ff184cdf", -- 57e0
		x"10014e75", -- 57e4
		x"48e7c088", -- 57e8
		x"42804281", -- 57ec
		x"2878fed4", -- 57f0
		x"302c0056", -- 57f4
		x"08ac0005", -- 57f8
		x"000a671e", -- 57fc
		x"41fa01b9", -- 5800
		x"6100fef2", -- 5804
		x"322c0056", -- 5808
		x"302c00bc", -- 580c
		x"55404eac", -- 5810
		x"003c703f", -- 5814
		x"4eac0036", -- 5818
		x"600c6100", -- 581c
		x"fefa41fa", -- 5820
		x"01846100", -- 5824
		x"fed04cdf", -- 5828
		x"11034e75", -- 582c
		x"48e7c088", -- 5830
		x"2878fed4", -- 5834
		x"08ac0007", -- 5838
		x"000a4280", -- 583c
		x"4281302c", -- 5840
		x"0046e248", -- 5844
		x"5240322c", -- 5848
		x"00564eac", -- 584c
		x"003c0c6c", -- 5850
		x"0020032c", -- 5854
		x"660a41fa", -- 5858
		x"00c64eba", -- 585c
		x"fe8e6042", -- 5860
		x"41fa00d6", -- 5864
		x"4ebafe84", -- 5868
		x"594f204f", -- 586c
		x"4240102c", -- 5870
		x"032c6100", -- 5874
		x"b1b81017", -- 5878
		x"4eac0036", -- 587c
		x"102f0001", -- 5880
		x"0c000020", -- 5884
		x"6604103c", -- 5888
		x"00304eac", -- 588c
		x"0036584f", -- 5890
		x"102c032d", -- 5894
		x"4eac0036", -- 5898
		x"70204eac", -- 589c
		x"00364eac", -- 58a0
		x"00364cdf", -- 58a4
		x"11034e75", -- 58a8
		x"52414d20", -- 58ac
		x"4641494c", -- 58b0
		x"45442041", -- 58b4
		x"424f5645", -- 58b8
		x"20464646", -- 58bc
		x"46433030", -- 58c0
		x"30005241", -- 58c4
		x"4d20474f", -- 58c8
		x"4e452041", -- 58cc
		x"424f5645", -- 58d0
		x"20464646", -- 58d4
		x"46433030", -- 58d8
		x"30002054", -- 58dc
		x"65737469", -- 58e0
		x"6e67204d", -- 58e4
		x"656d6f72", -- 58e8
		x"7900204c", -- 58ec
		x"6f616469", -- 58f0
		x"6e67204d", -- 58f4
		x"656d6f72", -- 58f8
		x"79002042", -- 58fc
		x"6f6f7469", -- 5900
		x"6e672053", -- 5904
		x"79737465", -- 5908
		x"6d002053", -- 590c
		x"79737465", -- 5910
		x"6d205365", -- 5914
		x"61726368", -- 5918
		x"204d6f64", -- 591c
		x"65002057", -- 5920
		x"61697469", -- 5924
		x"6e672053", -- 5928
		x"79737465", -- 592c
		x"6d205365", -- 5930
		x"6c656374", -- 5934
		x"696f6e00", -- 5938
		x"20537973", -- 593c
		x"74656d20", -- 5940
		x"53656c65", -- 5944
		x"63746564", -- 5948
		x"20697320", -- 594c
		x"00205365", -- 5950
		x"61726368", -- 5954
		x"20506175", -- 5958
		x"73656420", -- 595c
		x"28454e54", -- 5960
		x"45522054", -- 5964
		x"6f20436f", -- 5968
		x"6e74696e", -- 596c
		x"75652900", -- 5970
		x"20536561", -- 5974
		x"72636820", -- 5978
		x"50617573", -- 597c
		x"65642028", -- 5980
		x"52455455", -- 5984
		x"524e2054", -- 5988
		x"6f20436f", -- 598c
		x"6e74696e", -- 5990
		x"75652900", -- 5994
		x"2053656c", -- 5998
		x"662d5465", -- 599c
		x"7374204d", -- 59a0
		x"6f646500", -- 59a4
		x"20524553", -- 59a8
		x"45542054", -- 59ac
		x"6f20506f", -- 59b0
		x"7765722d", -- 59b4
		x"55700020", -- 59b8
		x"52455345", -- 59bc
		x"5420546f", -- 59c0
		x"20506f77", -- 59c4
		x"65722d55", -- 59c8
		x"702c2053", -- 59cc
		x"50414345", -- 59d0
		x"20636c65", -- 59d4
		x"61727320", -- 59d8
		x"696e7075", -- 59dc
		x"74002043", -- 59e0
		x"6f6e7469", -- 59e4
		x"6e756520", -- 59e8
		x"6174204f", -- 59ec
		x"776e2052", -- 59f0
		x"69736b20", -- 59f4
		x"28454e54", -- 59f8
		x"45522054", -- 59fc
		x"6f20436f", -- 5a00
		x"6e74696e", -- 5a04
		x"75652900", -- 5a08
		x"20436f6e", -- 5a0c
		x"74696e75", -- 5a10
		x"65206174", -- 5a14
		x"204f776e", -- 5a18
		x"20526973", -- 5a1c
		x"6b202852", -- 5a20
		x"45545552", -- 5a24
		x"4e20546f", -- 5a28
		x"20436f6e", -- 5a2c
		x"74696e75", -- 5a30
		x"65290020", -- 5a34
		x"57616974", -- 5a38
		x"696e6720", -- 5a3c
		x"31204d69", -- 5a40
		x"6e757465", -- 5a44
		x"2028454e", -- 5a48
		x"54455220", -- 5a4c
		x"746f2041", -- 5a50
		x"626f7274", -- 5a54
		x"20576169", -- 5a58
		x"74290020", -- 5a5c
		x"57616974", -- 5a60
		x"696e6720", -- 5a64
		x"31204d69", -- 5a68
		x"6e757465", -- 5a6c
		x"20285245", -- 5a70
		x"5455524e", -- 5a74
		x"20746f20", -- 5a78
		x"41626f72", -- 5a7c
		x"74205761", -- 5a80
		x"69742900", -- 5a84
		x"20554e45", -- 5a88
		x"58504543", -- 5a8c
		x"54454420", -- 5a90
		x"55534520", -- 5a94
		x"4f462000", -- 5a98
		x"204e4f54", -- 5a9c
		x"20454e4f", -- 5aa0
		x"55474820", -- 5aa4
		x"4d454d4f", -- 5aa8
		x"52590020", -- 5aac
		x"53595354", -- 5ab0
		x"454d2057", -- 5ab4
		x"4f554c44", -- 5ab8
		x"204c4f41", -- 5abc
		x"4420544f", -- 5ac0
		x"4f204849", -- 5ac4
		x"47480020", -- 5ac8
		x"53595354", -- 5acc
		x"454d204e", -- 5ad0
		x"4f542046", -- 5ad4
		x"4f554e44", -- 5ad8
		x"00436f70", -- 5adc
		x"79726967", -- 5ae0
		x"68742031", -- 5ae4
		x"3938392c", -- 5ae8
		x"00486577", -- 5aec
		x"6c657474", -- 5af0
		x"2d506163", -- 5af4
		x"6b617264", -- 5af8
		x"20436f6d", -- 5afc
		x"70616e79", -- 5b00
		x"2e00416c", -- 5b04
		x"6c205269", -- 5b08
		x"67687473", -- 5b0c
		x"20526573", -- 5b10
		x"65727665", -- 5b14
		x"642e0020", -- 5b18
		x"004d4336", -- 5b1c
		x"38303030", -- 5b20
		x"2050726f", -- 5b24
		x"63657373", -- 5b28
		x"6f720000", -- 5b2c
		x"416c7068", -- 5b30
		x"61205669", -- 5b34
		x"64656f00", -- 5b38
		x"42697420", -- 5b3c
		x"4d617070", -- 5b40
		x"65642056", -- 5b44
		x"6964656f", -- 5b48
		x"0048502d", -- 5b4c
		x"48494c2e", -- 5b50
		x"4b657962", -- 5b54
		x"6f617264", -- 5b58
		x"00436f6e", -- 5b5c
		x"736f6c65", -- 5b60
		x"204b6579", -- 5b64
		x"626f6172", -- 5b68
		x"64206174", -- 5b6c
		x"20202000", -- 5b70
		x"436f6c6f", -- 5b74
		x"72204772", -- 5b78
		x"61706869", -- 5b7c
		x"63730047", -- 5b80
		x"72617068", -- 5b84
		x"69637300", -- 5b88
		x"48502d49", -- 5b8c
		x"42004850", -- 5b90
		x"39383632", -- 5b94
		x"3000444d", -- 5b98
		x"412d0048", -- 5b9c
		x"50393836", -- 5ba0
		x"33350048", -- 5ba4
		x"50393832", -- 5ba8
		x"34380046", -- 5bac
		x"5020436f", -- 5bb0
		x"70726f63", -- 5bb4
		x"6573736f", -- 5bb8
		x"72004d43", -- 5bbc
		x"36383838", -- 5bc0
		x"3120436f", -- 5bc4
		x"70726f63", -- 5bc8
		x"6573736f", -- 5bcc
		x"72004d43", -- 5bd0
		x"36383838", -- 5bd4
		x"3220436f", -- 5bd8
		x"70726f63", -- 5bdc
		x"6573736f", -- 5be0
		x"72004850", -- 5be4
		x"39383238", -- 5be8
		x"3620436f", -- 5bec
		x"70726f63", -- 5bf0
		x"6573736f", -- 5bf4
		x"72002042", -- 5bf8
		x"79746573", -- 5bfc
		x"004d656d", -- 5c00
		x"6f727920", -- 5c04
		x"4661696c", -- 5c08
		x"65642061", -- 5c0c
		x"7420004d", -- 5c10
		x"656d6f72", -- 5c14
		x"7920476f", -- 5c18
		x"6e652061", -- 5c1c
		x"74200044", -- 5c20
		x"61746120", -- 5c24
		x"50617269", -- 5c28
		x"74792045", -- 5c2c
		x"72726f72", -- 5c30
		x"20617420", -- 5c34
		x"00506172", -- 5c38
		x"69747920", -- 5c3c
		x"42697420", -- 5c40
		x"4572726f", -- 5c44
		x"72206174", -- 5c48
		x"20002049", -- 5c4c
		x"676e6f72", -- 5c50
		x"65640020", -- 5c54
		x"61742000", -- 5c58
		x"20466169", -- 5c5c
		x"6c656400", -- 5c60
		x"20506173", -- 5c64
		x"73656400", -- 5c68
		x"53595354", -- 5c6c
		x"454d5f00", -- 5c70
		x"53595300", -- 5c74
		x"00000000", -- 5c78
		x"00005265", -- 5c7c
		x"6d6f7465", -- 5c80
		x"20436f6e", -- 5c84
		x"736f6c65", -- 5c88
		x"20617420", -- 5c8c
		x"00436f6e", -- 5c90
		x"66696775", -- 5c94
		x"72617469", -- 5c98
		x"6f6e2045", -- 5c9c
		x"4550524f", -- 5ca0
		x"4d200001", -- 5ca4
		x"48503938", -- 5ca8
		x"36323420", -- 5cac
		x"2848502d", -- 5cb0
		x"49422900", -- 5cb4
		x"02485039", -- 5cb8
		x"38363236", -- 5cbc
		x"20285253", -- 5cc0
		x"2d323332", -- 5cc4
		x"29004248", -- 5cc8
		x"50393836", -- 5ccc
		x"34342028", -- 5cd0
		x"52532d32", -- 5cd4
		x"33322900", -- 5cd8
		x"03485039", -- 5cdc
		x"38363232", -- 5ce0
		x"20284750", -- 5ce4
		x"494f2900", -- 5ce8
		x"04485039", -- 5cec
		x"38363233", -- 5cf0
		x"20284243", -- 5cf4
		x"44290005", -- 5cf8
		x"48503938", -- 5cfc
		x"36343220", -- 5d00
		x"2852532d", -- 5d04
		x"32333220", -- 5d08
		x"4d555829", -- 5d0c
		x"00064850", -- 5d10
		x"20504152", -- 5d14
		x"414c4c45", -- 5d18
		x"4c000748", -- 5d1c
		x"50393832", -- 5d20
		x"36352028", -- 5d24
		x"53435349", -- 5d28
		x"20532033", -- 5d2c
		x"32290027", -- 5d30
		x"48503938", -- 5d34
		x"32363520", -- 5d38
		x"28534353", -- 5d3c
		x"49205320", -- 5d40
		x"31362900", -- 5d44
		x"47485039", -- 5d48
		x"38323635", -- 5d4c
		x"20285343", -- 5d50
		x"53492044", -- 5d54
		x"20333229", -- 5d58
		x"00674850", -- 5d5c
		x"39383236", -- 5d60
		x"35202853", -- 5d64
		x"43534920", -- 5d68
		x"44203136", -- 5d6c
		x"29000848", -- 5d70
		x"50393836", -- 5d74
		x"32352028", -- 5d78
		x"48532048", -- 5d7c
		x"502d4942", -- 5d80
		x"29004848", -- 5d84
		x"502d4942", -- 5d88
		x"20284853", -- 5d8c
		x"20333229", -- 5d90
		x"00094850", -- 5d94
		x"2d48494c", -- 5d98
		x"2e4b6579", -- 5d9c
		x"626f6172", -- 5da0
		x"64000c48", -- 5da4
		x"50393836", -- 5da8
		x"34370011", -- 5dac
		x"48503938", -- 5db0
		x"36343620", -- 5db4
		x"28564d45", -- 5db8
		x"29003148", -- 5dbc
		x"50393835", -- 5dc0
		x"37372028", -- 5dc4
		x"564d4529", -- 5dc8
		x"00514850", -- 5dcc
		x"20453134", -- 5dd0
		x"38304120", -- 5dd4
		x"28565849", -- 5dd8
		x"29001248", -- 5ddc
		x"50393836", -- 5de0
		x"34300015", -- 5de4
		x"48503938", -- 5de8
		x"36343320", -- 5dec
		x"284c414e", -- 5df0
		x"29001648", -- 5df4
		x"50393836", -- 5df8
		x"39350019", -- 5dfc
		x"42697420", -- 5e00
		x"4d617070", -- 5e04
		x"65642056", -- 5e08
		x"6964656f", -- 5e0c
		x"00394269", -- 5e10
		x"74204d61", -- 5e14
		x"70706564", -- 5e18
		x"20566964", -- 5e1c
		x"656f001b", -- 5e20
		x"48503938", -- 5e24
		x"32353300", -- 5e28
		x"1c485039", -- 5e2c
		x"38363237", -- 5e30
		x"001d4850", -- 5e34
		x"39383633", -- 5e38
		x"33001e48", -- 5e3c
		x"50393832", -- 5e40
		x"35392028", -- 5e44
		x"42554229", -- 5e48
		x"00004944", -- 5e4c
		x"00485039", -- 5e50
		x"38363238", -- 5e54
		x"20285253", -- 5e58
		x"2d323332", -- 5e5c
		x"290048e7", -- 5e60
		x"80802078", -- 5e64
		x"fed46100", -- 5e68
		x"f6a40838", -- 5e6c
		x"0000fed2", -- 5e70
		x"6718317c", -- 5e74
		x"00320046", -- 5e78
		x"217c0051", -- 5e7c
		x"27040042", -- 5e80
		x"217c0051", -- 5e84
		x"2704004e", -- 5e88
		x"6016317c", -- 5e8c
		x"00500046", -- 5e90
		x"217c0051", -- 5e94
		x"21a00042", -- 5e98
		x"217c0051", -- 5e9c
		x"21a0004e", -- 5ea0
		x"31680046", -- 5ea4
		x"004ce3e8", -- 5ea8
		x"004c317c", -- 5eac
		x"00190056", -- 5eb0
		x"30280056", -- 5eb4
		x"c0e8004c", -- 5eb8
		x"d0a80042", -- 5ebc
		x"21400052", -- 5ec0
		x"317c4ef9", -- 5ec4
		x"0030217c", -- 5ec8
		x"00005e62", -- 5ecc
		x"0032317c", -- 5ed0
		x"4ef9003c", -- 5ed4
		x"217c0000", -- 5ed8
		x"6160003e", -- 5edc
		x"317c4ef9", -- 5ee0
		x"0036217c", -- 5ee4
		x"00006058", -- 5ee8
		x"00387001", -- 5eec
		x"6100f828", -- 5ef0
		x"2f3c000b", -- 5ef4
		x"71b04eba", -- 5ef8
		x"f3724cdf", -- 5efc
		x"01014e75", -- 5f00
		x"48e7f8f8", -- 5f04
		x"6100f3b4", -- 5f08
		x"6100f784", -- 5f0c
		x"2078fed4", -- 5f10
		x"610000ea", -- 5f14
		x"0c82ffff", -- 5f18
		x"ffff6608", -- 5f1c
		x"4cdf1f1f", -- 5f20
		x"600002e2", -- 5f24
		x"3142004c", -- 5f28
		x"2078fed4", -- 5f2c
		x"20680048", -- 5f30
		x"61000080", -- 5f34
		x"2078fed4", -- 5f38
		x"21430042", -- 5f3c
		x"24680048", -- 5f40
		x"224ad2c2", -- 5f44
		x"12290000", -- 5f48
		x"050a0011", -- 5f4c
		x"02820000", -- 5f50
		x"ffff0241", -- 5f54
		x"00ff84c1", -- 5f58
		x"31420056", -- 5f5c
		x"030a000d", -- 5f60
		x"10290002", -- 5f64
		x"02810000", -- 5f68
		x"ffff0240", -- 5f6c
		x"00ff82c0", -- 5f70
		x"31410046", -- 5f74
		x"217c0000", -- 5f78
		x"0000004e", -- 5f7c
		x"c4c12142", -- 5f80
		x"0052317c", -- 5f84
		x"4ef90030", -- 5f88
		x"217c0000", -- 5f8c
		x"5f040032", -- 5f90
		x"317c4ef9", -- 5f94
		x"003c217c", -- 5f98
		x"000061be", -- 5f9c
		x"003e317c", -- 5fa0
		x"4ef90036", -- 5fa4
		x"217c0000", -- 5fa8
		x"60820038", -- 5fac
		x"4cdf1f1f", -- 5fb0
		x"4e752f01", -- 5fb4
		x"12280001", -- 5fb8
		x"02010060", -- 5fbc
		x"672c4283", -- 5fc0
		x"42810308", -- 5fc4
		x"005d1630", -- 5fc8
		x"1800223c", -- 5fcc
		x"00000010", -- 5fd0
		x"e3abb1fc", -- 5fd4
		x"01000000", -- 5fd8
		x"6d02d688", -- 5fdc
		x"bffc0000", -- 5fe0
		x"01006304", -- 5fe4
		x"221f4e75", -- 5fe8
		x"4ed41628", -- 5fec
		x"4001c6bc", -- 5ff0
		x"0000000f", -- 5ff4
		x"223c0000", -- 5ff8
		x"001460d4", -- 5ffc
		x"48e740e0", -- 6000
		x"323cfffc", -- 6004
		x"2078fed4", -- 6008
		x"20680048", -- 600c
		x"42820508", -- 6010
		x"003b2248", -- 6014
		x"b47c0000", -- 6018
		x"672cd3c2", -- 601c
		x"42421429", -- 6020
		x"00004a02", -- 6024
		x"67205342", -- 6028
		x"5c410c31", -- 602c
		x"00011000", -- 6030
		x"670651ca", -- 6034
		x"fff4600e", -- 6038
		x"45f11002", -- 603c
		x"050a0000", -- 6040
		x"4cdf0702", -- 6044
		x"4e7508ec", -- 6048
		x"0004005c", -- 604c
		x"243cffff", -- 6050
		x"ffff60ec", -- 6054
		x"48e780c0", -- 6058
		x"2278fed4", -- 605c
		x"2069004e", -- 6060
		x"40e7007c", -- 6064
		x"070030c0", -- 6068
		x"b1e90052", -- 606c
		x"6d042069", -- 6070
		x"00422348", -- 6074
		x"004e46df", -- 6078
		x"4cdf0301", -- 607c
		x"4e7548e7", -- 6080
		x"fff02278", -- 6084
		x"fed42069", -- 6088
		x"004840e7", -- 608c
		x"007c0700", -- 6090
		x"42823429", -- 6094
		x"004c45f0", -- 6098
		x"28004241", -- 609c
		x"4242122a", -- 60a0
		x"0000142a", -- 60a4
		x"00022829", -- 60a8
		x"004e3629", -- 60ac
		x"004688c3", -- 60b0
		x"36044844", -- 60b4
		x"c8c20b08", -- 60b8
		x"0005c6c1", -- 60bc
		x"cac3da84", -- 60c0
		x"26690042", -- 60c4
		x"d7c52e0b", -- 60c8
		x"0c000020", -- 60cc
		x"66000022", -- 60d0
		x"0b080005", -- 60d4
		x"48c55342", -- 60d8
		x"53417800", -- 60dc
		x"360216c4", -- 60e0
		x"51cbfffc", -- 60e4
		x"de852647", -- 60e8
		x"51c9fff2", -- 60ec
		x"60000050", -- 60f0
		x"16025e03", -- 60f4
		x"e60be30b", -- 60f8
		x"024300ff", -- 60fc
		x"c6c1902a", -- 6100
		x"00060280", -- 6104
		x"000000ff", -- 6108
		x"c6c03c01", -- 610c
		x"53463002", -- 6110
		x"1832380a", -- 6114
		x"7a070b04", -- 6118
		x"56db5340", -- 611c
		x"670851cd", -- 6120
		x"fff65483", -- 6124
		x"60ea4a46", -- 6128
		x"67140b08", -- 612c
		x"00050285", -- 6130
		x"0000ffff", -- 6134
		x"de852647", -- 6138
		x"548351ce", -- 613c
		x"ffd252a9", -- 6140
		x"004e2029", -- 6144
		x"004eb0a9", -- 6148
		x"00526d08", -- 614c
		x"237c0000", -- 6150
		x"0000004e", -- 6154
		x"46df4cdf", -- 6158
		x"0fff4e75", -- 615c
		x"48e7f080", -- 6160
		x"40e7007c", -- 6164
		x"07002078", -- 6168
		x"fed42428", -- 616c
		x"004e94a8", -- 6170
		x"004284e8", -- 6174
		x"004c3602", -- 6178
		x"4842e24a", -- 617c
		x"4a006f0e", -- 6180
		x"488048c0", -- 6184
		x"538080e8", -- 6188
		x"00464840", -- 618c
		x"34004a01", -- 6190
		x"6f0e4881", -- 6194
		x"48c15381", -- 6198
		x"82e80056", -- 619c
		x"48413601", -- 61a0
		x"c6e8004c", -- 61a4
		x"d642d642", -- 61a8
		x"48c3d6a8", -- 61ac
		x"00422143", -- 61b0
		x"004e46df", -- 61b4
		x"4cdf010f", -- 61b8
		x"4e7548e7", -- 61bc
		x"e08040e7", -- 61c0
		x"007c0700", -- 61c4
		x"2078fed4", -- 61c8
		x"2428004e", -- 61cc
		x"84e80046", -- 61d0
		x"4a016604", -- 61d4
		x"12025201", -- 61d8
		x"4a006606", -- 61dc
		x"48421002", -- 61e0
		x"52005301", -- 61e4
		x"53000280", -- 61e8
		x"000000ff", -- 61ec
		x"02810000", -- 61f0
		x"00ffc2e8", -- 61f4
		x"0046d081", -- 61f8
		x"2140004e", -- 61fc
		x"46df4cdf", -- 6200
		x"01074e75", -- 6204
		x"2f082078", -- 6208
		x"fed4317c", -- 620c
		x"00500046", -- 6210
		x"317c0019", -- 6214
		x"0056317c", -- 6218
		x"4ef90030", -- 621c
		x"217c0000", -- 6220
		x"62080032", -- 6224
		x"317c4ef9", -- 6228
		x"003c217c", -- 622c
		x"00006246", -- 6230
		x"003e317c", -- 6234
		x"4ef90036", -- 6238
		x"217c0000", -- 623c
		x"62460038", -- 6240
		x"205f4e75", -- 6244
		x"302dfffe", -- 6248
		x"2078fed4", -- 624c
		x"2228005e", -- 6250
		x"41f8fdd2", -- 6254
		x"610000ca", -- 6258
		x"421841f8", -- 625c
		x"fdd26100", -- 6260
		x"f51c41f8", -- 6264
		x"fdd230fc", -- 6268
		x"2020610a", -- 626c
		x"421841f8", -- 6270
		x"fdd26000", -- 6274
		x"f50848e7", -- 6278
		x"e0400c00", -- 627c
		x"00026610", -- 6280
		x"0281e200", -- 6284
		x"00000c81", -- 6288
		x"e2000000", -- 628c
		x"66027008", -- 6290
		x"43fa002a", -- 6294
		x"1419670a", -- 6298
		x"b0026706", -- 629c
		x"4a1966fc", -- 62a0
		x"60f210d9", -- 62a4
		x"66fc117c", -- 62a8
		x"0020ffff", -- 62ac
		x"b07c0008", -- 62b0
		x"63046100", -- 62b4
		x"a7984cdf", -- 62b8
		x"02074e75", -- 62bc
		x"014e6f20", -- 62c0
		x"44657669", -- 62c4
		x"63650002", -- 62c8
		x"4e6f204d", -- 62cc
		x"65646975", -- 62d0
		x"6d00034e", -- 62d4
		x"6f742052", -- 62d8
		x"65616479", -- 62dc
		x"00045265", -- 62e0
		x"61642045", -- 62e4
		x"72726f72", -- 62e8
		x"00054261", -- 62ec
		x"64204861", -- 62f0
		x"72647761", -- 62f4
		x"72650006", -- 62f8
		x"42616420", -- 62fc
		x"53746174", -- 6300
		x"65000742", -- 6304
		x"75732045", -- 6308
		x"72726f72", -- 630c
		x"00084e6f", -- 6310
		x"20536572", -- 6314
		x"76657200", -- 6318
		x"00457272", -- 631c
		x"6f720000", -- 6320
		x"48e7ff78", -- 6324
		x"10fc003a", -- 6328
		x"48e740c0", -- 632c
		x"2278fed4", -- 6330
		x"2f29005e", -- 6334
		x"2341005e", -- 6338
		x"598f2f08", -- 633c
		x"6100ee6e", -- 6340
		x"245f1412", -- 6344
		x"2078fed4", -- 6348
		x"215f005e", -- 634c
		x"4cdf0302", -- 6350
		x"24484240", -- 6354
		x"101a5340", -- 6358
		x"6d0410da", -- 635c
		x"60f80802", -- 6360
		x"00036708", -- 6364
		x"10fc002c", -- 6368
		x"10fc0020", -- 636c
		x"e0990802", -- 6370
		x"00006708", -- 6374
		x"42401001", -- 6378
		x"6100a6d2", -- 637c
		x"08020004", -- 6380
		x"670810fc", -- 6384
		x"002c10fc", -- 6388
		x"00200802", -- 638c
		x"00066732", -- 6390
		x"2278fed4", -- 6394
		x"45e90000", -- 6398
		x"2248201a", -- 639c
		x"6100e718", -- 63a0
		x"30126100", -- 63a4
		x"e7202049", -- 63a8
		x"2278fed4", -- 63ac
		x"10fc0020", -- 63b0
		x"45e900ce", -- 63b4
		x"4240101a", -- 63b8
		x"660210da", -- 63bc
		x"51c8fffc", -- 63c0
		x"6050e199", -- 63c4
		x"42401001", -- 63c8
		x"08020001", -- 63cc
		x"67100802", -- 63d0
		x"00046706", -- 63d4
		x"6100a676", -- 63d8
		x"60046100", -- 63dc
		x"a69ce199", -- 63e0
		x"e1990802", -- 63e4
		x"0002672a", -- 63e8
		x"10fc002c", -- 63ec
		x"10fc0020", -- 63f0
		x"42401001", -- 63f4
		x"08020005", -- 63f8
		x"6714c07c", -- 63fc
		x"000f6100", -- 6400
		x"a64c1001", -- 6404
		x"e84810fc", -- 6408
		x"002c10fc", -- 640c
		x"00206100", -- 6410
		x"a63c4cdf", -- 6414
		x"1eff4e75", -- 6418
		x"48e70070", -- 641c
		x"2278fed4", -- 6420
		x"246900aa", -- 6424
		x"266900ae", -- 6428
		x"2f2f000c", -- 642c
		x"4e7561e8", -- 6430
		x"61000042", -- 6434
		x"4cdf0e00", -- 6438
		x"584f4e75", -- 643c
		x"61da6100", -- 6440
		x"00584cdf", -- 6444
		x"0e00584f", -- 6448
		x"4e7561cc", -- 644c
		x"610000a6", -- 6450
		x"4cdf0e00", -- 6454
		x"584f4e75", -- 6458
		x"61be6100", -- 645c
		x"00a04cdf", -- 6460
		x"0e00584f", -- 6464
		x"4e7561b0", -- 6468
		x"6100009a", -- 646c
		x"4cdf0e00", -- 6470
		x"584f4e75", -- 6474
		x"48e70060", -- 6478
		x"2278fed4", -- 647c
		x"246900aa", -- 6480
		x"08120000", -- 6484
		x"66fa4cdf", -- 6488
		x"06004e75", -- 648c
		x"44fc0000", -- 6490
		x"4e7544fc", -- 6494
		x"00044e75", -- 6498
		x"4a806750", -- 649c
		x"08380001", -- 64a0
		x"feda663c", -- 64a4
		x"80fc00c8", -- 64a8
		x"02800000", -- 64ac
		x"ffff0640", -- 64b0
		x"00012f00", -- 64b4
		x"48576100", -- 64b8
		x"ed38201f", -- 64bc
		x"90bc0000", -- 64c0
		x"00092f00", -- 64c4
		x"48574eba", -- 64c8
		x"ed52201f", -- 64cc
		x"08120001", -- 64d0
		x"67be2f00", -- 64d4
		x"48574eba", -- 64d8
		x"ed626aee", -- 64dc
		x"588f7000", -- 64e0
		x"08120001", -- 64e4
		x"57c8fffa", -- 64e8
		x"66a24e75", -- 64ec
		x"08120001", -- 64f0
		x"66fa4e75", -- 64f4
		x"61a26698", -- 64f8
		x"14816096", -- 64fc
		x"619a6690", -- 6500
		x"1681608e", -- 6504
		x"4a80675c", -- 6508
		x"08380001", -- 650c
		x"feda663e", -- 6510
		x"80fc00c8", -- 6514
		x"02800000", -- 6518
		x"ffff0640", -- 651c
		x"00012f00", -- 6520
		x"48576100", -- 6524
		x"eccc201f", -- 6528
		x"90bc0000", -- 652c
		x"00092f00", -- 6530
		x"48574eba", -- 6534
		x"ece6201f", -- 6538
		x"08120000", -- 653c
		x"6600001c", -- 6540
		x"2f004857", -- 6544
		x"4ebaecf4", -- 6548
		x"6aec588f", -- 654c
		x"70000812", -- 6550
		x"000056c8", -- 6554
		x"fffa6700", -- 6558
		x"ff344280", -- 655c
		x"12121013", -- 6560
		x"6000ff30", -- 6564
		x"08120000", -- 6568
		x"66f060f8", -- 656c
		x"428148e7", -- 6570
		x"00702278", -- 6574
		x"fed42469", -- 6578
		x"00aa2669", -- 657c
		x"00ae6184", -- 6580
		x"4cdf0e00", -- 6584
		x"6600ff0a", -- 6588
		x"08810000", -- 658c
		x"08010007", -- 6590
		x"6700fefe", -- 6594
		x"08010006", -- 6598
		x"665a0c00", -- 659c
		x"003c6d00", -- 65a0
		x"fef02400", -- 65a4
		x"4840943c", -- 65a8
		x"003c08c1", -- 65ac
		x"00000801", -- 65b0
		x"00046606", -- 65b4
		x"d4bc0000", -- 65b8
		x"00422078", -- 65bc
		x"fed44a28", -- 65c0
		x"00a9671c", -- 65c4
		x"2f031628", -- 65c8
		x"00a84883", -- 65cc
		x"e54b207c", -- 65d0
		x"0000680c", -- 65d4
		x"20703000", -- 65d8
		x"10302800", -- 65dc
		x"261f6006", -- 65e0
		x"2042103b", -- 65e4
		x"80140801", -- 65e8
		x"00056604", -- 65ec
		x"0200001f", -- 65f0
		x"48404e75", -- 65f4
		x"72004e75", -- 65f8
		x"302e2c2b", -- 65fc
		x"3132332d", -- 6600
		x"3435362a", -- 6604
		x"3738392f", -- 6608
		x"4528295e", -- 660c
		x"31323334", -- 6610
		x"35363738", -- 6614
		x"39302d3d", -- 6618
		x"5b5d3b27", -- 661c
		x"2c2e2f20", -- 6620
		x"4f504b4c", -- 6624
		x"51574552", -- 6628
		x"54595549", -- 662c
		x"41534446", -- 6630
		x"47484a4d", -- 6634
		x"5a584356", -- 6638
		x"424e7f60", -- 663c
		x"7cf1b0b3", -- 6640
		x"df7eebef", -- 6644
		x"f5f0f6f7", -- 6648
		x"fa5cd1f4", -- 664c
		x"fbd12140", -- 6650
		x"2324255e", -- 6654
		x"262a2829", -- 6658
		x"5f2b7b7d", -- 665c
		x"3a223c3e", -- 6660
		x"3f206f70", -- 6664
		x"6b6c7177", -- 6668
		x"65727479", -- 666c
		x"75696173", -- 6670
		x"64666768", -- 6674
		x"6a6d7a78", -- 6678
		x"6376626e", -- 667c
		x"302e2c2b", -- 6680
		x"3132332d", -- 6684
		x"3435362a", -- 6688
		x"3738392f", -- 668c
		x"4528295e", -- 6690
		x"31323334", -- 6694
		x"35363738", -- 6698
		x"39302d3d", -- 669c
		x"5b5d3b27", -- 66a0
		x"2c2e2f20", -- 66a4
		x"4f504b4c", -- 66a8
		x"51574552", -- 66ac
		x"545a5549", -- 66b0
		x"41534446", -- 66b4
		x"47484a4d", -- 66b8
		x"59584356", -- 66bc
		x"424e302e", -- 66c0
		x"2c2b3132", -- 66c4
		x"332d3435", -- 66c8
		x"362a3738", -- 66cc
		x"392f4528", -- 66d0
		x"295e2140", -- 66d4
		x"2324255e", -- 66d8
		x"262a2829", -- 66dc
		x"5f2b7b7d", -- 66e0
		x"3a343c3e", -- 66e4
		x"3f206f70", -- 66e8
		x"6b6c7177", -- 66ec
		x"6572747a", -- 66f0
		x"75696173", -- 66f4
		x"64666768", -- 66f8
		x"6a6d7978", -- 66fc
		x"6376626e", -- 6700
		x"302e2c2b", -- 6704
		x"3132332d", -- 6708
		x"3435362a", -- 670c
		x"3738392f", -- 6710
		x"4528295e", -- 6714
		x"21402324", -- 6718
		x"255e262a", -- 671c
		x"28292d3d", -- 6720
		x"5b5d4d27", -- 6724
		x"2c2e2f20", -- 6728
		x"4f504b4c", -- 672c
		x"515a4552", -- 6730
		x"54595549", -- 6734
		x"41534446", -- 6738
		x"47484a2c", -- 673c
		x"57584356", -- 6740
		x"424e302e", -- 6744
		x"2c2b3132", -- 6748
		x"332d3435", -- 674c
		x"362a3738", -- 6750
		x"392f4528", -- 6754
		x"295e3132", -- 6758
		x"33343536", -- 675c
		x"37383930", -- 6760
		x"5f2b7b7d", -- 6764
		x"6d343c3e", -- 6768
		x"3f206f70", -- 676c
		x"6b6c717a", -- 6770
		x"65727479", -- 6774
		x"75696173", -- 6778
		x"64666768", -- 677c
		x"6a3f7778", -- 6780
		x"6376626e", -- 6784
		x"302e2c2b", -- 6788
		x"3132332d", -- 678c
		x"3435362a", -- 6790
		x"3738392f", -- 6794
		x"4528295e", -- 6798
		x"21402324", -- 679c
		x"255e262a", -- 67a0
		x"28292d3d", -- 67a4
		x"5b5d4d27", -- 67a8
		x"2c2e2f20", -- 67ac
		x"4f504b4c", -- 67b0
		x"415a4552", -- 67b4
		x"54595549", -- 67b8
		x"51534446", -- 67bc
		x"47484a2c", -- 67c0
		x"57584356", -- 67c4
		x"424e302e", -- 67c8
		x"2c2b3132", -- 67cc
		x"332d3435", -- 67d0
		x"362a3738", -- 67d4
		x"392f4528", -- 67d8
		x"295e3132", -- 67dc
		x"33343536", -- 67e0
		x"37383930", -- 67e4
		x"5f2b7b7d", -- 67e8
		x"6d343c3e", -- 67ec
		x"3f206f70", -- 67f0
		x"6b6c617a", -- 67f4
		x"65727479", -- 67f8
		x"75697173", -- 67fc
		x"64666768", -- 6800
		x"6a3f7778", -- 6804
		x"6376626e", -- 6808
		x"000065fc", -- 680c
		x"000065fc", -- 6810
		x"000065fc", -- 6814
		x"00006680", -- 6818
		x"000065fc", -- 681c
		x"000065fc", -- 6820
		x"000065fc", -- 6824
		x"000065fc", -- 6828
		x"000065fc", -- 682c
		x"000065fc", -- 6830
		x"000065fc", -- 6834
		x"00006704", -- 6838
		x"000065fc", -- 683c
		x"000065fc", -- 6840
		x"000065fc", -- 6844
		x"00006680", -- 6848
		x"000065fc", -- 684c
		x"000065fc", -- 6850
		x"000065fc", -- 6854
		x"000065fc", -- 6858
		x"000065fc", -- 685c
		x"00006788", -- 6860
		x"000065fc", -- 6864
		x"000065fc", -- 6868
		x"000065fc", -- 686c
		x"00006680", -- 6870
		x"000065fc", -- 6874
		x"00006788", -- 6878
		x"000065fc", -- 687c
		x"000065fc", -- 6880
		x"000065fc", -- 6884
		x"000065fc", -- 6888
		x"48e7e070", -- 688c
		x"2278fed4", -- 6890
		x"246900aa", -- 6894
		x"266900ae", -- 6898
		x"428072a3", -- 689c
		x"6100fc56", -- 68a0
		x"32026100", -- 68a4
		x"fc58e049", -- 68a8
		x"6100fc52", -- 68ac
		x"4cdf0e07", -- 68b0
		x"4e750838", -- 68b4
		x"0003fed2", -- 68b8
		x"661e0c2c", -- 68bc
		x"00ff00a6", -- 68c0
		x"6716343c", -- 68c4
		x"08f861c0", -- 68c8
		x"2f3c0004", -- 68cc
		x"93e04eba", -- 68d0
		x"e99a343c", -- 68d4
		x"08f861b0", -- 68d8
		x"4e7548e7", -- 68dc
		x"00602278", -- 68e0
		x"fed42469", -- 68e4
		x"00aa14bc", -- 68e8
		x"00b20838", -- 68ec
		x"0003fed2", -- 68f0
		x"66100839", -- 68f4
		x"00020047", -- 68f8
		x"800566f6", -- 68fc
		x"4cdf0600", -- 6900
		x"4e732469", -- 6904
		x"00b20812", -- 6908
		x"000366fa", -- 690c
		x"60ee48e7", -- 6910
		x"e0702278", -- 6914
		x"fed42469", -- 6918
		x"00aa2669", -- 691c
		x"00ae4280", -- 6920
		x"1412725f", -- 6924
		x"6100fbce", -- 6928
		x"72b26100", -- 692c
		x"fbc86100", -- 6930
		x"fbc46100", -- 6934
		x"fb64613c", -- 6938
		x"613a0801", -- 693c
		x"00014cdf", -- 6940
		x"0e07660c", -- 6944
		x"48790088", -- 6948
		x"00244eba", -- 694c
		x"e2ca584f", -- 6950
		x"2f0c2878", -- 6954
		x"fed4082c", -- 6958
		x"0001005c", -- 695c
		x"670a197c", -- 6960
		x"0002005d", -- 6964
		x"285f4e73", -- 6968
		x"1c38fed2", -- 696c
		x"41fa9a8e", -- 6970
		x"6000da48", -- 6974
		x"6100fb76", -- 6978
		x"14bc0005", -- 697c
		x"10120800", -- 6980
		x"000166f8", -- 6984
		x"08000000", -- 6988
		x"67f21213", -- 698c
		x"c07c00f0", -- 6990
		x"b07c0040", -- 6994
		x"66e64e75", -- 6998
		x"48e780f0", -- 699c
		x"2278fed4", -- 69a0
		x"48e72006", -- 69a4
		x"45f90060", -- 69a8
		x"00004242", -- 69ac
		x"b47c0020", -- 69b0
		x"6c000044", -- 69b4
		x"4dfa0034", -- 69b8
		x"2a4f701f", -- 69bc
		x"c02a0001", -- 69c0
		x"0c400009", -- 69c4
		x"6700008a", -- 69c8
		x"b03c001c", -- 69cc
		x"6714b03c", -- 69d0
		x"001d670e", -- 69d4
		x"b03c001a", -- 69d8
		x"66105442", -- 69dc
		x"d5fc0002", -- 69e0
		x"00005242", -- 69e4
		x"d5fc0001", -- 69e8
		x"00005242", -- 69ec
		x"d5fc0001", -- 69f0
		x"00002e4d", -- 69f4
		x"60b64cdf", -- 69f8
		x"600442a9", -- 69fc
		x"00b240e7", -- 6a00
		x"337c4ef9", -- 6a04
		x"0300237c", -- 6a08
		x"0000699c", -- 6a0c
		x"03026000", -- 6a10
		x"016a2e4d", -- 6a14
		x"08e90005", -- 6a18
		x"005c41fa", -- 6a1c
		x"f13d6100", -- 6a20
		x"e4606100", -- 6a24
		x"000460ce", -- 6a28
		x"48e7fee0", -- 6a2c
		x"72007015", -- 6a30
		x"4ea9003c", -- 6a34
		x"43f8fdd2", -- 6a38
		x"300248c0", -- 6a3c
		x"6100e048", -- 6a40
		x"421141f8", -- 6a44
		x"fdd26100", -- 6a48
		x"eca24cdf", -- 6a4c
		x"077f4e75", -- 6a50
		x"70236100", -- 6a54
		x"e3dc4dfa", -- 6a58
		x"ffba4a2a", -- 6a5c
		x"0003234a", -- 6a60
		x"00b2264a", -- 6a64
		x"d5fc0000", -- 6a68
		x"500cd7fc", -- 6a6c
		x"00005004", -- 6a70
		x"234a00aa", -- 6a74
		x"234b00ae", -- 6a78
		x"203c0007", -- 6a7c
		x"a1206100", -- 6a80
		x"fa84668e", -- 6a84
		x"c23c00f0", -- 6a88
		x"0c010070", -- 6a8c
		x"66840c00", -- 6a90
		x"008e6600", -- 6a94
		x"ff7e41fa", -- 6a98
		x"f0c16100", -- 6a9c
		x"e3e06188", -- 6aa0
		x"4cdf6004", -- 6aa4
		x"602448e7", -- 6aa8
		x"80f02278", -- 6aac
		x"fed4247c", -- 6ab0
		x"00428003", -- 6ab4
		x"234a00aa", -- 6ab8
		x"267c0042", -- 6abc
		x"8001234b", -- 6ac0
		x"00ae237c", -- 6ac4
		x"00420000", -- 6ac8
		x"00b240e7", -- 6acc
		x"007c0700", -- 6ad0
		x"10121013", -- 6ad4
		x"70a06100", -- 6ad8
		x"010e4200", -- 6adc
		x"61000100", -- 6ae0
		x"610000fc", -- 6ae4
		x"610000f8", -- 6ae8
		x"70016100", -- 6aec
		x"00f2705c", -- 6af0
		x"610000f4", -- 6af4
		x"422900a9", -- 6af8
		x"70116100", -- 6afc
		x"00ea6100", -- 6b00
		x"00ee0800", -- 6b04
		x"00056710", -- 6b08
		x"02000007", -- 6b0c
		x"0c000002", -- 6b10
		x"6706137c", -- 6b14
		x"000100a9", -- 6b18
		x"70126100", -- 6b1c
		x"00ca6100", -- 6b20
		x"00ce1340", -- 6b24
		x"00a80c29", -- 6b28
		x"000100a9", -- 6b2c
		x"6614303c", -- 6b30
		x"0000323c", -- 6b34
		x"00eb4eba", -- 6b38
		x"f9bc323c", -- 6b3c
		x"00974eba", -- 6b40
		x"f9bc31fc", -- 6b44
		x"4ef9ffbe", -- 6b48
		x"21fc0000", -- 6b4c
		x"6c56ffc0", -- 6b50
		x"31fc4ef9", -- 6b54
		x"ff3421fc", -- 6b58
		x"00006912", -- 6b5c
		x"ff3631fc", -- 6b60
		x"4ef9ff9a", -- 6b64
		x"21fc0000", -- 6b68
		x"4d20ff9c", -- 6b6c
		x"337c4ef9", -- 6b70
		x"0300237c", -- 6b74
		x"00006aaa", -- 6b78
		x"0302337c", -- 6b7c
		x"4ef90306", -- 6b80
		x"237c0000", -- 6b84
		x"6c0e0308", -- 6b88
		x"337c4ef9", -- 6b8c
		x"030c237c", -- 6b90
		x"00006c22", -- 6b94
		x"030e08a9", -- 6b98
		x"0003000b", -- 6b9c
		x"42690322", -- 6ba0
		x"337c0312", -- 6ba4
		x"0324337c", -- 6ba8
		x"03120326", -- 6bac
		x"4229032c", -- 6bb0
		x"137c0020", -- 6bb4
		x"032d6100", -- 6bb8
		x"08d46100", -- 6bbc
		x"09340838", -- 6bc0
		x"0003fed2", -- 6bc4
		x"67104aa9", -- 6bc8
		x"00b2670a", -- 6bcc
		x"246900b2", -- 6bd0
		x"08ea0007", -- 6bd4
		x"000346df", -- 6bd8
		x"4cdf0f01", -- 6bdc
		x"4e756100", -- 6be0
		x"f90c1680", -- 6be4
		x"4e756100", -- 6be8
		x"f9041480", -- 6bec
		x"4e751012", -- 6bf0
		x"08000000", -- 6bf4
		x"67f81f13", -- 6bf8
		x"c07c00f0", -- 6bfc
		x"b03c0040", -- 6c00
		x"6704101f", -- 6c04
		x"60e8101f", -- 6c08
		x"4e752f08", -- 6c0c
		x"2078fed4", -- 6c10
		x"4a680322", -- 6c14
		x"670444fc", -- 6c18
		x"0000205f", -- 6c1c
		x"4e7548e7", -- 6c20
		x"40c02278", -- 6c24
		x"fed44ea9", -- 6c28
		x"030667fa", -- 6c2c
		x"32290324", -- 6c30
		x"41f11000", -- 6c34
		x"10105269", -- 6c38
		x"03245369", -- 6c3c
		x"03220c69", -- 6c40
		x"03220324", -- 6c44
		x"6606337c", -- 6c48
		x"03120324", -- 6c4c
		x"4cdf0302", -- 6c50
		x"4e7548e7", -- 6c54
		x"e0c02278", -- 6c58
		x"fed44280", -- 6c5c
		x"48e70030", -- 6c60
		x"246900aa", -- 6c64
		x"266900ae", -- 6c68
		x"12121013", -- 6c6c
		x"4cdf0c00", -- 6c70
		x"08010007", -- 6c74
		x"670000f8", -- 6c78
		x"08010006", -- 6c7c
		x"660000f0", -- 6c80
		x"08e90003", -- 6c84
		x"000b0801", -- 6c88
		x"00056700", -- 6c8c
		x"00dc0c40", -- 6c90
		x"002e6606", -- 6c94
		x"70086000", -- 6c98
		x"00900c40", -- 6c9c
		x"00396606", -- 6ca0
		x"700d6000", -- 6ca4
		x"00840c00", -- 6ca8
		x"003c6d00", -- 6cac
		x"00bc0c00", -- 6cb0
		x"007d6e00", -- 6cb4
		x"00b46100", -- 6cb8
		x"f8ea4840", -- 6cbc
		x"08e90003", -- 6cc0
		x"000b0c29", -- 6cc4
		x"000000a9", -- 6cc8
		x"66260c29", -- 6ccc
		x"000200a8", -- 6cd0
		x"661eb03c", -- 6cd4
		x"00596712", -- 6cd8
		x"b03c005a", -- 6cdc
		x"670cb03c", -- 6ce0
		x"00796706", -- 6ce4
		x"b03c007a", -- 6ce8
		x"66060a00", -- 6cec
		x"00036038", -- 6cf0
		x"b03c0020", -- 6cf4
		x"6732b03c", -- 6cf8
		x"000d672c", -- 6cfc
		x"b03c0008", -- 6d00
		x"6726b03c", -- 6d04
		x"00306548", -- 6d08
		x"b03c0039", -- 6d0c
		x"631ab03c", -- 6d10
		x"0041653c", -- 6d14
		x"b03c005a", -- 6d18
		x"630eb03c", -- 6d1c
		x"00616530", -- 6d20
		x"b03c007a", -- 6d24
		x"63026028", -- 6d28
		x"0c690010", -- 6d2c
		x"03226720", -- 6d30
		x"32290326", -- 6d34
		x"41f11000", -- 6d38
		x"10805269", -- 6d3c
		x"03260c69", -- 6d40
		x"03220326", -- 6d44
		x"6606337c", -- 6d48
		x"03120326", -- 6d4c
		x"52690322", -- 6d50
		x"08290007", -- 6d54
		x"00a6660e", -- 6d58
		x"4a29004c", -- 6d5c
		x"670808e9", -- 6d60
		x"0000004d", -- 6d64
		x"6008610c", -- 6d68
		x"226900c2", -- 6d6c
		x"4e914cdf", -- 6d70
		x"03074e73", -- 6d74
		x"48e7e0c0", -- 6d78
		x"40e7007c", -- 6d7c
		x"07002278", -- 6d80
		x"fed408e9", -- 6d84
		x"000600c0", -- 6d88
		x"72001229", -- 6d8c
		x"00ba7400", -- 6d90
		x"142900bb", -- 6d94
		x"206900b6", -- 6d98
		x"08290007", -- 6d9c
		x"00c06700", -- 6da0
		x"009a08a9", -- 6da4
		x"000300c0", -- 6da8
		x"67046100", -- 6dac
		x"00f408a9", -- 6db0
		x"000400c0", -- 6db4
		x"670c4ea9", -- 6db8
		x"03066778", -- 6dbc
		x"4ea9030c", -- 6dc0
		x"60f40c01", -- 6dc4
		x"0000676c", -- 6dc8
		x"b4016508", -- 6dcc
		x"08290000", -- 6dd0
		x"00c06760", -- 6dd4
		x"4ea90306", -- 6dd8
		x"67604ea9", -- 6ddc
		x"030cb03c", -- 6de0
		x"000d6614", -- 6de4
		x"08290000", -- 6de8
		x"00c06648", -- 6dec
		x"11801000", -- 6df0
		x"08e90001", -- 6df4
		x"00c0603c", -- 6df8
		x"b03c0008", -- 6dfc
		x"66104a02", -- 6e00
		x"67d25302", -- 6e04
		x"11bc0020", -- 6e08
		x"20006140", -- 6e0c
		x"60c6b03c", -- 6e10
		x"001f63c0", -- 6e14
		x"b03c0020", -- 6e18
		x"660c0829", -- 6e1c
		x"000200c0", -- 6e20
		x"6704617c", -- 6e24
		x"60aeb401", -- 6e28
		x"64a21180", -- 6e2c
		x"2000611c", -- 6e30
		x"52026094", -- 6e34
		x"08a90007", -- 6e38
		x"00c01342", -- 6e3c
		x"00bb08a9", -- 6e40
		x"000600c0", -- 6e44
		x"46df4cdf", -- 6e48
		x"03074e75", -- 6e4c
		x"48e7d800", -- 6e50
		x"302900bc", -- 6e54
		x"322900be", -- 6e58
		x"36023829", -- 6e5c
		x"00465744", -- 6e60
		x"b0446610", -- 6e64
		x"b2690056", -- 6e68
		x"660a2f29", -- 6e6c
		x"004e7600", -- 6e70
		x"50c46004", -- 6e74
		x"d04251c4", -- 6e78
		x"4ea9003c", -- 6e7c
		x"10303000", -- 6e80
		x"4ea90036", -- 6e84
		x"5243b642", -- 6e88
		x"63f24a44", -- 6e8c
		x"670c235f", -- 6e90
		x"004e7000", -- 6e94
		x"72004ea9", -- 6e98
		x"003c4cdf", -- 6e9c
		x"001b4e75", -- 6ea0
		x"48e7c800", -- 6ea4
		x"2f29004e", -- 6ea8
		x"302900bc", -- 6eac
		x"322900be", -- 6eb0
		x"4ea9003c", -- 6eb4
		x"70206008", -- 6eb8
		x"11802110", -- 6ebc
		x"4ea90036", -- 6ec0
		x"51cafff6", -- 6ec4
		x"74003029", -- 6ec8
		x"00bc3229", -- 6ecc
		x"00be3829", -- 6ed0
		x"00465744", -- 6ed4
		x"b044660e", -- 6ed8
		x"b2690056", -- 6edc
		x"66082357", -- 6ee0
		x"004e7000", -- 6ee4
		x"72004ea9", -- 6ee8
		x"003c588f", -- 6eec
		x"4cdf0013", -- 6ef0
		x"4e752f0c", -- 6ef4
		x"2878fed4", -- 6ef8
		x"422c005d", -- 6efc
		x"08ec0001", -- 6f00
		x"005c285f", -- 6f04
		x"4e752f09", -- 6f08
		x"40e7007c", -- 6f0c
		x"07002278", -- 6f10
		x"fed408a9", -- 6f14
		x"0001005c", -- 6f18
		x"4a29005d", -- 6f1c
		x"671a0c29", -- 6f20
		x"0002005d", -- 6f24
		x"67062269", -- 6f28
		x"00c24e91", -- 6f2c
		x"1c38fed2", -- 6f30
		x"41fa94ca", -- 6f34
		x"6000d484", -- 6f38
		x"46df225f", -- 6f3c
		x"4e755228", -- 6f40
		x"004c6100", -- 6f44
		x"fe305328", -- 6f48
		x"004c6608", -- 6f4c
		x"08a80000", -- 6f50
		x"004d66ea", -- 6f54
		x"4e752f08", -- 6f58
		x"2078fed4", -- 6f5c
		x"317c0050", -- 6f60
		x"0046317c", -- 6f64
		x"00180056", -- 6f68
		x"317c0000", -- 6f6c
		x"0058317c", -- 6f70
		x"0002005a", -- 6f74
		x"317c0001", -- 6f78
		x"004e317c", -- 6f7c
		x"00180050", -- 6f80
		x"2168004e", -- 6f84
		x"00524228", -- 6f88
		x"004c4228", -- 6f8c
		x"004d317c", -- 6f90
		x"4ef90030", -- 6f94
		x"217c0000", -- 6f98
		x"6f5a0032", -- 6f9c
		x"317c4ef9", -- 6fa0
		x"003c217c", -- 6fa4
		x"00007086", -- 6fa8
		x"003e317c", -- 6fac
		x"4ef90036", -- 6fb0
		x"217c0000", -- 6fb4
		x"6fd40038", -- 6fb8
		x"5228004c", -- 6fbc
		x"40e7007c", -- 6fc0
		x"07006100", -- 6fc4
		x"015a46df", -- 6fc8
		x"6100ff7c", -- 6fcc
		x"205f4e75", -- 6fd0
		x"48e7f080", -- 6fd4
		x"2078fed4", -- 6fd8
		x"5228004c", -- 6fdc
		x"40e7007c", -- 6fe0
		x"07003228", -- 6fe4
		x"00583428", -- 6fe8
		x"00520c00", -- 6fec
		x"00206616", -- 6ff0
		x"08280006", -- 6ff4
		x"00c0665e", -- 6ff8
		x"3601d642", -- 6ffc
		x"b6680046", -- 7000
		x"6c745241", -- 7004
		x"606c0c00", -- 7008
		x"001f622e", -- 700c
		x"0c00000d", -- 7010
		x"66067400", -- 7014
		x"7200603e", -- 7018
		x"0c00000a", -- 701c
		x"66085268", -- 7020
		x"00545342", -- 7024
		x"60300c00", -- 7028
		x"0008664a", -- 702c
		x"53416e42", -- 7030
		x"72005542", -- 7034
		x"6e207401", -- 7038
		x"602e4840", -- 703c
		x"303c0020", -- 7040
		x"60066100", -- 7044
		x"03605242", -- 7048
		x"51c9fff8", -- 704c
		x"72004840", -- 7050
		x"317c0002", -- 7054
		x"005a6100", -- 7058
		x"034c5242", -- 705c
		x"b4680046", -- 7060
		x"6f067401", -- 7064
		x"52680054", -- 7068
		x"31420052", -- 706c
		x"21680052", -- 7070
		x"004e3141", -- 7074
		x"005846df", -- 7078
		x"6100fecc", -- 707c
		x"4cdf010f", -- 7080
		x"4e7548e7", -- 7084
		x"f8802078", -- 7088
		x"fed45228", -- 708c
		x"004c40e7", -- 7090
		x"007c0700", -- 7094
		x"317c0000", -- 7098
		x"00583428", -- 709c
		x"00523828", -- 70a0
		x"00465744", -- 70a4
		x"b0446d06", -- 70a8
		x"b2680056", -- 70ac
		x"671e4a41", -- 70b0
		x"66043228", -- 70b4
		x"00503628", -- 70b8
		x"00549641", -- 70bc
		x"67063141", -- 70c0
		x"0054615a", -- 70c4
		x"4a406604", -- 70c8
		x"3028004e", -- 70cc
		x"34280052", -- 70d0
		x"31400052", -- 70d4
		x"3600b443", -- 70d8
		x"672e6e0e", -- 70dc
		x"70206100", -- 70e0
		x"02c45242", -- 70e4
		x"b4436df4", -- 70e8
		x"601e5744", -- 70ec
		x"b4446c0c", -- 70f0
		x"70086100", -- 70f4
		x"02b07020", -- 70f8
		x"610002aa", -- 70fc
		x"70086100", -- 7100
		x"02a45342", -- 7104
		x"b4436ee4", -- 7108
		x"31420052", -- 710c
		x"21680052", -- 7110
		x"004e46df", -- 7114
		x"6100fe30", -- 7118
		x"4cdf011f", -- 711c
		x"4e7548e7", -- 7120
		x"80802078", -- 7124
		x"fed44a68", -- 7128
		x"005a6f1c", -- 712c
		x"700d6100", -- 7130
		x"0274700a", -- 7134
		x"6100026e", -- 7138
		x"317c0001", -- 713c
		x"0052317c", -- 7140
		x"00000058", -- 7144
		x"5368005a", -- 7148
		x"4cdf0101", -- 714c
		x"4e7548e7", -- 7150
		x"ffce0838", -- 7154
		x"0001fed9", -- 7158
		x"6600018e", -- 715c
		x"2878fed4", -- 7160
		x"207c0060", -- 7164
		x"00004dfa", -- 7168
		x"01522a4f", -- 716c
		x"74001428", -- 7170
		x"00010882", -- 7174
		x"00076700", -- 7178
		x"01460c02", -- 717c
		x"00026710", -- 7180
		x"0c020005", -- 7184
		x"67000062", -- 7188
		x"0c020042", -- 718c
		x"66000130", -- 7190
		x"52886100", -- 7194
		x"d8445388", -- 7198
		x"4a006600", -- 719c
		x"01227043", -- 71a0
		x"0c020042", -- 71a4
		x"67041028", -- 71a8
		x"0007ec08", -- 71ac
		x"194000a6", -- 71b0
		x"294800a2", -- 71b4
		x"43f8fdd2", -- 71b8
		x"41faeac0", -- 71bc
		x"12d866fc", -- 71c0
		x"5349701f", -- 71c4
		x"c06c00a2", -- 71c8
		x"6100d8bc", -- 71cc
		x"421941f8", -- 71d0
		x"fdd26100", -- 71d4
		x"e5a8397c", -- 71d8
		x"0001032e", -- 71dc
		x"61000110", -- 71e0
		x"6100fd74", -- 71e4
		x"60000102", -- 71e8
		x"48e700a0", -- 71ec
		x"24486100", -- 71f0
		x"001c4cdf", -- 71f4
		x"05004a00", -- 71f8
		x"67046000", -- 71fc
		x"00c2d1fc", -- 7200
		x"00004000", -- 7204
		x"197c0004", -- 7208
		x"00a660a4", -- 720c
		x"4dfa007c", -- 7210
		x"40c1d5fc", -- 7214
		x"00004000", -- 7218
		x"203c0000", -- 721c
		x"0bb80838", -- 7220
		x"0001feda", -- 7224
		x"66422f3c", -- 7228
		x"000001f4", -- 722c
		x"48574eba", -- 7230
		x"dfc04857", -- 7234
		x"4ebadfe4", -- 7238
		x"201f41fa", -- 723c
		x"fffe007c", -- 7240
		x"0700082a", -- 7244
		x"0007c005", -- 7248
		x"6600006c", -- 724c
		x"082a0004", -- 7250
		x"4001663a", -- 7254
		x"422ac005", -- 7258
		x"46c12f00", -- 725c
		x"48574eba", -- 7260
		x"dfda6ad4", -- 7264
		x"588f7000", -- 7268
		x"41fafffe", -- 726c
		x"007c0700", -- 7270
		x"082a0007", -- 7274
		x"c005663e", -- 7278
		x"082a0004", -- 727c
		x"4001660e", -- 7280
		x"422ac005", -- 7284
		x"46c151c8", -- 7288
		x"ffe050c0", -- 728c
		x"4e7508aa", -- 7290
		x"00044001", -- 7294
		x"422ac005", -- 7298
		x"46c10c2a", -- 729c
		x"00e04e47", -- 72a0
		x"67100c2a", -- 72a4
		x"000d4e47", -- 72a8
		x"67080c2a", -- 72ac
		x"000c4e47", -- 72b0
		x"66d84200", -- 72b4
		x"4e7546c1", -- 72b8
		x"4ed02e4d", -- 72bc
		x"74000202", -- 72c0
		x"001f7004", -- 72c4
		x"0c02001a", -- 72c8
		x"67107002", -- 72cc
		x"0c02001c", -- 72d0
		x"67080c02", -- 72d4
		x"001d6702", -- 72d8
		x"70014840", -- 72dc
		x"d1c0b1fc", -- 72e0
		x"00800000", -- 72e4
		x"6500fe80", -- 72e8
		x"4cdf73ff", -- 72ec
		x"4e7548e7", -- 72f0
		x"e0c82878", -- 72f4
		x"fed4206c", -- 72f8
		x"00a20c2c", -- 72fc
		x"008000a6", -- 7300
		x"67000054", -- 7304
		x"0c2c0004", -- 7308
		x"00a66750", -- 730c
		x"707cc02c", -- 7310
		x"00a66642", -- 7314
		x"707fc028", -- 7318
		x"0001720e", -- 731c
		x"74430c00", -- 7320
		x"00426708", -- 7324
		x"12280005", -- 7328
		x"14280007", -- 732c
		x"c27c000f", -- 7330
		x"e34943fb", -- 7334
		x"1050117c", -- 7338
		x"00800017", -- 733c
		x"11590013", -- 7340
		x"11510011", -- 7344
		x"c43c003f", -- 7348
		x"11420017", -- 734c
		x"117c0005", -- 7350
		x"001351ec", -- 7354
		x"00a74cdf", -- 7358
		x"13074e75", -- 735c
		x"7430720f", -- 7360
		x"11424e25", -- 7364
		x"11414e27", -- 7368
		x"143c0001", -- 736c
		x"610003c8", -- 7370
		x"51ec00a7", -- 7374
		x"08280007", -- 7378
		x"c00366da", -- 737c
		x"08e80007", -- 7380
		x"c00360d2", -- 7384
		x"0c000800", -- 7388
		x"05740476", -- 738c
		x"04000300", -- 7390
		x"02000100", -- 7394
		x"00800055", -- 7398
		x"0040002b", -- 739c
		x"00200015", -- 73a0
		x"00100008", -- 73a4
		x"48e7f088", -- 73a8
		x"2878fed4", -- 73ac
		x"206c00a2", -- 73b0
		x"7200122c", -- 73b4
		x"00a6b27c", -- 73b8
		x"00046700", -- 73bc
		x"0088647e", -- 73c0
		x"e341323b", -- 73c4
		x"10064efb", -- 73c8
		x"1002003e", -- 73cc
		x"005e0066", -- 73d0
		x"00660828", -- 73d4
		x"00060003", -- 73d8
		x"660c4e75", -- 73dc
		x"08280006", -- 73e0
		x"c0036602", -- 73e4
		x"4e750838", -- 73e8
		x"0004feda", -- 73ec
		x"67104267", -- 73f0
		x"487affe8", -- 73f4
		x"40e7007c", -- 73f8
		x"07006000", -- 73fc
		x"016e0838", -- 7400
		x"0002feda", -- 7404
		x"67e860e8", -- 7408
		x"532c00a7", -- 740c
		x"6a2261c2", -- 7410
		x"08280005", -- 7414
		x"001b67f6", -- 7418
		x"117c0005", -- 741c
		x"001161b2", -- 7420
		x"4a2c00a7", -- 7424
		x"6a0a60f6", -- 7428
		x"61a84a2c", -- 742c
		x"00a766f8", -- 7430
		x"61a00828", -- 7434
		x"0005001b", -- 7438
		x"67f61140", -- 743c
		x"00114cdf", -- 7440
		x"110f4e75", -- 7444
		x"61964a2c", -- 7448
		x"00a766f8", -- 744c
		x"618e4242", -- 7450
		x"14284e1b", -- 7454
		x"16021202", -- 7458
		x"d43c000e", -- 745c
		x"0202000f", -- 7460
		x"b4284e13", -- 7464
		x"67e61401", -- 7468
		x"d44249e8", -- 746c
		x"4f211980", -- 7470
		x"20005241", -- 7474
		x"0201000f", -- 7478
		x"11414e1b", -- 747c
		x"b6284e13", -- 7480
		x"66bc143c", -- 7484
		x"00026100", -- 7488
		x"02ae60b2", -- 748c
		x"48e78088", -- 7490
		x"2878fed4", -- 7494
		x"206c00a2", -- 7498
		x"0c2c0004", -- 749c
		x"00a6671e", -- 74a0
		x"707cc02c", -- 74a4
		x"00a66610", -- 74a8
		x"08280005", -- 74ac
		x"001b67f8", -- 74b0
		x"08280006", -- 74b4
		x"001b67f0", -- 74b8
		x"4cdf1101", -- 74bc
		x"4e751028", -- 74c0
		x"4e1bb028", -- 74c4
		x"4e1366f6", -- 74c8
		x"6100ff08", -- 74cc
		x"60ea48e7", -- 74d0
		x"808840e7", -- 74d4
		x"007c0700", -- 74d8
		x"10284e13", -- 74dc
		x"b0284e1b", -- 74e0
		x"670a5240", -- 74e4
		x"0200000f", -- 74e8
		x"11404e1b", -- 74ec
		x"46df60c8", -- 74f0
		x"48e7e088", -- 74f4
		x"2878fed4", -- 74f8
		x"206c00a2", -- 74fc
		x"4a2c00a6", -- 7500
		x"6b366100", -- 7504
		x"fdea7030", -- 7508
		x"0c2c0004", -- 750c
		x"00a6672e", -- 7510
		x"727cc22c", -- 7514
		x"00a66620", -- 7518
		x"117c0080", -- 751c
		x"0003c028", -- 7520
		x"0003e848", -- 7524
		x"c0fc0006", -- 7528
		x"41f8ffb2", -- 752c
		x"90c030fc", -- 7530
		x"4ef920fc", -- 7534
		x"0000756e", -- 7538
		x"4cdf1107", -- 753c
		x"4e75323c", -- 7540
		x"0100343c", -- 7544
		x"000249e8", -- 7548
		x"4c0118c2", -- 754c
		x"528c51c9", -- 7550
		x"fffa6100", -- 7554
		x"ff7ac028", -- 7558
		x"c0030828", -- 755c
		x"0007c003", -- 7560
		x"66c008e8", -- 7564
		x"0007c003", -- 7568
		x"60b848e7", -- 756c
		x"e0c02278", -- 7570
		x"fed42069", -- 7574
		x"00a20c29", -- 7578
		x"000400a6", -- 757c
		x"670000a4", -- 7580
		x"10280015", -- 7584
		x"0c000004", -- 7588
		x"672e0828", -- 758c
		x"00070003", -- 7590
		x"67160828", -- 7594
		x"0004001b", -- 7598
		x"670e0829", -- 759c
		x"0001005c", -- 75a0
		x"670a137c", -- 75a4
		x"0002005d", -- 75a8
		x"6000f7c4", -- 75ac
		x"1c38fed2", -- 75b0
		x"41fa8e4a", -- 75b4
		x"6000ce04", -- 75b8
		x"10280011", -- 75bc
		x"72001229", -- 75c0
		x"00a6b27c", -- 75c4
		x"000464e0", -- 75c8
		x"e341323b", -- 75cc
		x"10064efb", -- 75d0
		x"10020008", -- 75d4
		x"0016002e", -- 75d8
		x"002e0c00", -- 75dc
		x"00066620", -- 75e0
		x"137c004e", -- 75e4
		x"00a760c0", -- 75e8
		x"0c000011", -- 75ec
		x"660651e9", -- 75f0
		x"00a760b4", -- 75f4
		x"0c000013", -- 75f8
		x"660650e9", -- 75fc
		x"00a760a8", -- 7600
		x"08280007", -- 7604
		x"000367a0", -- 7608
		x"6000f6b2", -- 760c
		x"42284e41", -- 7610
		x"4e714228", -- 7614
		x"40014e71", -- 7618
		x"4228c005", -- 761c
		x"4e7146df", -- 7620
		x"608640e7", -- 7624
		x"007c0700", -- 7628
		x"08280007", -- 762c
		x"c00566f8", -- 7630
		x"2f3c0000", -- 7634
		x"00324eba", -- 7638
		x"dc320828", -- 763c
		x"00014001", -- 7640
		x"67ca0828", -- 7644
		x"00014e41", -- 7648
		x"67c24228", -- 764c
		x"4e414e71", -- 7650
		x"42284001", -- 7654
		x"4e714228", -- 7658
		x"c0054e71", -- 765c
		x"46df7200", -- 7660
		x"12284e03", -- 7664
		x"1401d241", -- 7668
		x"48e71030", -- 766c
		x"47e84801", -- 7670
		x"b4284e0b", -- 7674
		x"66084cdf", -- 7678
		x"0c086000", -- 767c
		x"f6dc1033", -- 7680
		x"10005441", -- 7684
		x"16331000", -- 7688
		x"54415442", -- 768c
		x"024200ff", -- 7690
		x"024101ff", -- 7694
		x"11424e03", -- 7698
		x"08030004", -- 769c
		x"67084cdf", -- 76a0
		x"0c086000", -- 76a4
		x"fef60c00", -- 76a8
		x"00116606", -- 76ac
		x"51e900a7", -- 76b0
		x"60be0c00", -- 76b4
		x"00136606", -- 76b8
		x"50e900a7", -- 76bc
		x"60b20828", -- 76c0
		x"0007c003", -- 76c4
		x"67aa08e9", -- 76c8
		x"0003000b", -- 76cc
		x"b03c0020", -- 76d0
		x"6736b03c", -- 76d4
		x"000d6730", -- 76d8
		x"b03c0008", -- 76dc
		x"672ab03c", -- 76e0
		x"0030658c", -- 76e4
		x"b03c0039", -- 76e8
		x"631eb03c", -- 76ec
		x"00416580", -- 76f0
		x"b03c005a", -- 76f4
		x"6312b03c", -- 76f8
		x"00616500", -- 76fc
		x"ff74b03c", -- 7700
		x"007a6304", -- 7704
		x"6000ff6a", -- 7708
		x"0c690010", -- 770c
		x"03226700", -- 7710
		x"ff603229", -- 7714
		x"032645f1", -- 7718
		x"10001480", -- 771c
		x"52690326", -- 7720
		x"0c690322", -- 7724
		x"03266606", -- 7728
		x"337c0312", -- 772c
		x"03265269", -- 7730
		x"03226000", -- 7734
		x"ff3c40e7", -- 7738
		x"007c0700", -- 773c
		x"08280007", -- 7740
		x"c0056612", -- 7744
		x"85284e39", -- 7748
		x"00280002", -- 774c
		x"40034228", -- 7750
		x"c00546df", -- 7754
		x"4e7546d7", -- 7758
		x"60de48e7", -- 775c
		x"818e2878", -- 7760
		x"fed4207c", -- 7764
		x"00600000", -- 7768
		x"2e3c0002", -- 776c
		x"00002c7c", -- 7770
		x"0000779c", -- 7774
		x"2a4f1028", -- 7778
		x"00010c00", -- 777c
		x"001c671e", -- 7780
		x"d1c70200", -- 7784
		x"001f0c00", -- 7788
		x"001a6602", -- 778c
		x"d1c7b1fc", -- 7790
		x"00800000", -- 7794
		x"65d8602e", -- 7798
		x"2e4d4280", -- 779c
		x"60e248e7", -- 77a0
		x"00886100", -- 77a4
		x"d2944cdf", -- 77a8
		x"11004a00", -- 77ac
		x"66d22948", -- 77b0
		x"00a2d1fc", -- 77b4
		x"00010000", -- 77b8
		x"29480042", -- 77bc
		x"197c0080", -- 77c0
		x"00a66100", -- 77c4
		x"00984cdf", -- 77c8
		x"71814e75", -- 77cc
		x"48e7c0c0", -- 77d0
		x"2278fed4", -- 77d4
		x"20690042", -- 77d8
		x"91fc0000", -- 77dc
		x"80004280", -- 77e0
		x"323c17ff", -- 77e4
		x"20c020c0", -- 77e8
		x"20c020c0", -- 77ec
		x"51c9fff6", -- 77f0
		x"206900a2", -- 77f4
		x"117c0080", -- 77f8
		x"00014cdf", -- 77fc
		x"03034e75", -- 7800
		x"48e7c0c0", -- 7804
		x"2278fed4", -- 7808
		x"206900a2", -- 780c
		x"1029000b", -- 7810
		x"43fa002e", -- 7814
		x"08000000", -- 7818
		x"670443fa", -- 781c
		x"00324280", -- 7820
		x"720d1140", -- 7824
		x"00101159", -- 7828
		x"00125240", -- 782c
		x"51c9fff4", -- 7830
		x"4cdf0303", -- 7834
		x"4e7548e7", -- 7838
		x"c0c02278", -- 783c
		x"fed460cc", -- 7840
		x"29202203", -- 7844
		x"32053131", -- 7848
		x"00070000", -- 784c
		x"00002920", -- 7850
		x"22033d05", -- 7854
		x"31370007", -- 7858
		x"00000000", -- 785c
		x"6100ff6e", -- 7860
		x"2f0c2878", -- 7864
		x"fed4397c", -- 7868
		x"4ef90030", -- 786c
		x"297c0000", -- 7870
		x"78600032", -- 7874
		x"397c4ef9", -- 7878
		x"003c297c", -- 787c
		x"000061be", -- 7880
		x"003e397c", -- 7884
		x"4ef90036", -- 7888
		x"297c0000", -- 788c
		x"78b60038", -- 7890
		x"42ac004e", -- 7894
		x"397c0049", -- 7898
		x"0046397c", -- 789c
		x"00180056", -- 78a0
		x"297c0000", -- 78a4
		x"06d80052", -- 78a8
		x"08b80000", -- 78ac
		x"fed2285f", -- 78b0
		x"4e7548e7", -- 78b4
		x"f62840c6", -- 78b8
		x"007c2700", -- 78bc
		x"2878fed4", -- 78c0
		x"242c004e", -- 78c4
		x"22025241", -- 78c8
		x"b26c0052", -- 78cc
		x"66024281", -- 78d0
		x"2941004e", -- 78d4
		x"84ec0046", -- 78d8
		x"32024842", -- 78dc
		x"c2fc0380", -- 78e0
		x"c4fc0007", -- 78e4
		x"2602e68a", -- 78e8
		x"d282286c", -- 78ec
		x"0042d9c1", -- 78f0
		x"02430007", -- 78f4
		x"143b3056", -- 78f8
		x"4842143b", -- 78fc
		x"3048247c", -- 7900
		x"00002000", -- 7904
		x"024000ff", -- 7908
		x"e948d4c0", -- 790c
		x"303c000d", -- 7910
		x"4241121a", -- 7914
		x"e3094a03", -- 7918
		x"6702e679", -- 791c
		x"1a14ca02", -- 7920
		x"8a0118c5", -- 7924
		x"4842e059", -- 7928
		x"1a14ca02", -- 792c
		x"8a011885", -- 7930
		x"4842d9fc", -- 7934
		x"0000003f", -- 7938
		x"51c8ffd6", -- 793c
		x"46c64cdf", -- 7940
		x"146f4e75", -- 7944
		x"0180c0e0", -- 7948
		x"f0f8fcfe", -- 794c
		x"ffff7f3f", -- 7950
		x"1f0f0703", -- 7954
		x"60000026", -- 7958
		x"60000022", -- 795c
		x"6000001e", -- 7960
		x"600002ae", -- 7964
		x"600002a8", -- 7968
		x"600002a8", -- 796c
		x"6000000e", -- 7970
		x"6000029c", -- 7974
		x"60000298", -- 7978
		x"60000294", -- 797c
		x"3b7c0820", -- 7980
		x"fffe2e6d", -- 7984
		x"fff64e75", -- 7988
		x"42863c00", -- 798c
		x"2e068cfc", -- 7990
		x"03e84846", -- 7994
		x"42803006", -- 7998
		x"2f066100", -- 799c
		x"d0ea2c1f", -- 79a0
		x"12fc002c", -- 79a4
		x"48464280", -- 79a8
		x"30066100", -- 79ac
		x"d0da12fc", -- 79b0
		x"002041fa", -- 79b4
		x"0022be50", -- 79b8
		x"670c4a50", -- 79bc
		x"66044219", -- 79c0
		x"4e755888", -- 79c4
		x"60f03068", -- 79c8
		x"0002d1fc", -- 79cc
		x"000079da", -- 79d0
		x"6100d116", -- 79d4
		x"4e75042a", -- 79d8
		x"00740812", -- 79dc
		x"00910bfa", -- 79e0
		x"00ad0fe2", -- 79e4
		x"00bf0438", -- 79e8
		x"00d00820", -- 79ec
		x"00d00c08", -- 79f0
		x"00d01f90", -- 79f4
		x"00e52378", -- 79f8
		x"00e50439", -- 79fc
		x"00f30821", -- 7a00
		x"00f30c09", -- 7a04
		x"010b0ff1", -- 7a08
		x"011e13d9", -- 7a0c
		x"013017c1", -- 7a10
		x"01431ba9", -- 7a14
		x"0155043b", -- 7a18
		x"01700823", -- 7a1c
		x"0170043c", -- 7a20
		x"01800824", -- 7a24
		x"01990c0c", -- 7a28
		x"00f3043f", -- 7a2c
		x"01b30440", -- 7a30
		x"01cd17ca", -- 7a34
		x"01df1bb2", -- 7a38
		x"01df1f9a", -- 7a3c
		x"01f42382", -- 7a40
		x"020d2b52", -- 7a44
		x"02230000", -- 7a48
		x"0000494e", -- 7a4c
		x"4954202e", -- 7a50
		x"2e204241", -- 7a54
		x"44205452", -- 7a58
		x"41434b20", -- 7a5c
		x"30202c20", -- 7a60
		x"53494445", -- 7a64
		x"20300049", -- 7a68
		x"4e495420", -- 7a6c
		x"2e2e2054", -- 7a70
		x"4f4f204d", -- 7a74
		x"414e5920", -- 7a78
		x"42414420", -- 7a7c
		x"54524143", -- 7a80
		x"4b530049", -- 7a84
		x"4e495420", -- 7a88
		x"2e2e204c", -- 7a8c
		x"4f535420", -- 7a90
		x"44415441", -- 7a94
		x"00494e49", -- 7a98
		x"54202e2e", -- 7a9c
		x"2054494d", -- 7aa0
		x"45204f55", -- 7aa4
		x"5400444f", -- 7aa8
		x"4f52204f", -- 7aac
		x"50454e20", -- 7ab0
		x"2f204e4f", -- 7ab4
		x"204d4544", -- 7ab8
		x"4941004d", -- 7abc
		x"45444941", -- 7ac0
		x"20434841", -- 7ac4
		x"4e474544", -- 7ac8
		x"00534545", -- 7acc
		x"4b202e2e", -- 7ad0
		x"20545241", -- 7ad4
		x"434b204e", -- 7ad8
		x"4f542046", -- 7adc
		x"4f554e44", -- 7ae0
		x"00534545", -- 7ae4
		x"4b202e2e", -- 7ae8
		x"204e4f20", -- 7aec
		x"54524143", -- 7af0
		x"4b203000", -- 7af4
		x"52454144", -- 7af8
		x"202e2e20", -- 7afc
		x"4c4f5354", -- 7b00
		x"20444154", -- 7b04
		x"41005752", -- 7b08
		x"49544520", -- 7b0c
		x"2e2e204c", -- 7b10
		x"4f535420", -- 7b14
		x"44415441", -- 7b18
		x"00534545", -- 7b1c
		x"4b202e2e", -- 7b20
		x"204c4f53", -- 7b24
		x"54204441", -- 7b28
		x"54410057", -- 7b2c
		x"52495445", -- 7b30
		x"202e2e20", -- 7b34
		x"41444452", -- 7b38
		x"45535320", -- 7b3c
		x"43524320", -- 7b40
		x"4552524f", -- 7b44
		x"52004d45", -- 7b48
		x"44494120", -- 7b4c
		x"50524f54", -- 7b50
		x"45435445", -- 7b54
		x"44005245", -- 7b58
		x"4144202e", -- 7b5c
		x"2e205345", -- 7b60
		x"43544f52", -- 7b64
		x"204e4f54", -- 7b68
		x"20464f55", -- 7b6c
		x"4e440057", -- 7b70
		x"52495445", -- 7b74
		x"202e2e20", -- 7b78
		x"53454354", -- 7b7c
		x"4f52204e", -- 7b80
		x"4f542046", -- 7b84
		x"4f554e44", -- 7b88
		x"00534545", -- 7b8c
		x"4b202e2e", -- 7b90
		x"20414444", -- 7b94
		x"52455353", -- 7b98
		x"20435243", -- 7b9c
		x"20455252", -- 7ba0
		x"4f520052", -- 7ba4
		x"45414420", -- 7ba8
		x"2e2e2043", -- 7bac
		x"52432045", -- 7bb0
		x"52524f52", -- 7bb4
		x"00554e45", -- 7bb8
		x"58504543", -- 7bbc
		x"54454420", -- 7bc0
		x"494e5445", -- 7bc4
		x"52525550", -- 7bc8
		x"54005449", -- 7bcc
		x"4d454f55", -- 7bd0
		x"54204455", -- 7bd4
		x"52494e47", -- 7bd8
		x"20494e54", -- 7bdc
		x"45525255", -- 7be0
		x"50540049", -- 7be4
		x"4e544552", -- 7be8
		x"52555054", -- 7bec
		x"53204c4f", -- 7bf0
		x"434b4544", -- 7bf4
		x"204f5554", -- 7bf8
		x"00445249", -- 7bfc
		x"5645204e", -- 7c00
		x"4f542052", -- 7c04
		x"4553504f", -- 7c08
		x"4e44494e", -- 7c0c
		x"47004e75", -- 7c10
		x"4e730838", -- 7c14
		x"0001feda", -- 7c18
		x"662a48c0", -- 7c1c
		x"2f006700", -- 7c20
		x"00204857", -- 7c24
		x"4ebad5ca", -- 7c28
		x"48574eba", -- 7c2c
		x"d5ee0896", -- 7c30
		x"0002660c", -- 7c34
		x"48574eba", -- 7c38
		x"d6026af2", -- 7c3c
		x"08960002", -- 7c40
		x"588f4e75", -- 7c44
		x"223c0000", -- 7c48
		x"00c80896", -- 7c4c
		x"00026608", -- 7c50
		x"53816ef6", -- 7c54
		x"53406eec", -- 7c58
		x"4e7541fa", -- 7c5c
		x"d60e2948", -- 7c60
		x"036c41fa", -- 7c64
		x"d5b62948", -- 7c68
		x"037041fa", -- 7c6c
		x"d5e82948", -- 7c70
		x"037442ac", -- 7c74
		x"036442ac", -- 7c78
		x"036842ac", -- 7c7c
		x"037842ac", -- 7c80
		x"037c4280", -- 7c84
		x"102c00a9", -- 7c88
		x"39400354", -- 7c8c
		x"102c00a8", -- 7c90
		x"39400356", -- 7c94
		x"082c0004", -- 7c98
		x"000b6722", -- 7c9c
		x"4aac0010", -- 7ca0
		x"66044eba", -- 7ca4
		x"d1622038", -- 7ca8
		x"fdce2940", -- 7cac
		x"0380d0bc", -- 7cb0
		x"00000190", -- 7cb4
		x"29400384", -- 7cb8
		x"21c0fdce", -- 7cbc
		x"4e75204c", -- 7cc0
		x"91fc0001", -- 7cc4
		x"08002948", -- 7cc8
		x"0380d1fc", -- 7ccc
		x"00000190", -- 7cd0
		x"29480384", -- 7cd4
		x"4e752e42", -- 7cd8
		x"4cdf7fff", -- 7cdc
		x"4e7548e7", -- 7ce0
		x"fffe240f", -- 7ce4
		x"4dfafff0", -- 7ce8
		x"08b80005", -- 7cec
		x"fdcc47ec", -- 7cf0
		x"0340294a", -- 7cf4
		x"03444280", -- 7cf8
		x"010a0085", -- 7cfc
		x"4a8067d6", -- 7d00
		x"4bf20800", -- 7d04
		x"4a1566ce", -- 7d08
		x"4bed0004", -- 7d0c
		x"4a15671c", -- 7d10
		x"4a2d0002", -- 7d14
		x"66c04280", -- 7d18
		x"010d0004", -- 7d1c
		x"08000000", -- 7d20
		x"66b4e388", -- 7d24
		x"67b04bf5", -- 7d28
		x"080460e0", -- 7d2c
		x"4280010d", -- 7d30
		x"00040800", -- 7d34
		x"0000669e", -- 7d38
		x"2e00206c", -- 7d3c
		x"038443f0", -- 7d40
		x"08002949", -- 7d44
		x"03584bed", -- 7d48
		x"0008e288", -- 7d4c
		x"660c6086", -- 7d50
		x"090d0000", -- 7d54
		x"4bed0004", -- 7d58
		x"30c451c8", -- 7d5c
		x"fff448e7", -- 7d60
		x"ff80206c", -- 7d64
		x"03842807", -- 7d68
		x"4ebad13c", -- 7d6c
		x"4a404cdf", -- 7d70
		x"01ff6600", -- 7d74
		x"ff62294a", -- 7d78
		x"03447e02", -- 7d7c
		x"082c0000", -- 7d80
		x"000a6716", -- 7d84
		x"08380006", -- 7d88
		x"fed2660c", -- 7d8c
		x"08380007", -- 7d90
		x"fdcc6604", -- 7d94
		x"7e016002", -- 7d98
		x"7e032947", -- 7d9c
		x"0348296c", -- 7da0
		x"0380034c", -- 7da4
		x"297c0000", -- 7da8
		x"00000340", -- 7dac
		x"6118672c", -- 7db0
		x"bebc0000", -- 7db4
		x"00026700", -- 7db8
		x"ff1ebebc", -- 7dbc
		x"00000001", -- 7dc0
		x"67d67e02", -- 7dc4
		x"60d448e7", -- 7dc8
		x"fffe2f0b", -- 7dcc
		x"2a6c0384", -- 7dd0
		x"4e954cdf", -- 7dd4
		x"7fff4aac", -- 7dd8
		x"03604e75", -- 7ddc
		x"4dfa01ca", -- 7de0
		x"226c0380", -- 7de4
		x"4e55fff2", -- 7de8
		x"426dfff2", -- 7dec
		x"2b51fffc", -- 7df0
		x"0c070002", -- 7df4
		x"67562019", -- 7df8
		x"6f0001ae", -- 7dfc
		x"42863c2c", -- 7e00
		x"00565d46", -- 7e04
		x"bc806d00", -- 7e08
		x"01a0b0ad", -- 7e0c
		x"fffc6f04", -- 7e10
		x"2b40fffc", -- 7e14
		x"2b40fff4", -- 7e18
		x"29470348", -- 7e1c
		x"29400350", -- 7e20
		x"41f8fdd2", -- 7e24
		x"2948034c", -- 7e28
		x"197c0002", -- 7e2c
		x"03436196", -- 7e30
		x"66000176", -- 7e34
		x"2a2c035c", -- 7e38
		x"42305000", -- 7e3c
		x"61000202", -- 7e40
		x"20196cfc", -- 7e44
		x"0c80ffff", -- 7e48
		x"ffff67aa", -- 7e4c
		x"202dfffc", -- 7e50
		x"54802b40", -- 7e54
		x"fff8226c", -- 7e58
		x"03802b59", -- 7e5c
		x"fff42019", -- 7e60
		x"6c345989", -- 7e64
		x"0c070002", -- 7e68
		x"671841fa", -- 7e6c
		x"ddf44a6d", -- 7e70
		x"fff26706", -- 7e74
		x"6d0841fa", -- 7e78
		x"dde06100", -- 7e7c
		x"01f66100", -- 7e80
		x"02860c99", -- 7e84
		x"ffffffff", -- 7e88
		x"6600011e", -- 7e8c
		x"2b59fff4", -- 7e90
		x"426dfff2", -- 7e94
		x"60c8197c", -- 7e98
		x"00010343", -- 7e9c
		x"29400348", -- 7ea0
		x"6100ff24", -- 7ea4
		x"2c2c0360", -- 7ea8
		x"6f1c0c86", -- 7eac
		x"00000002", -- 7eb0
		x"67140c86", -- 7eb4
		x"00000003", -- 7eb8
		x"670c0c86", -- 7ebc
		x"00000006", -- 7ec0
		x"67046000", -- 7ec4
		x"00e442ac", -- 7ec8
		x"034841f8", -- 7ecc
		x"fdd22948", -- 7ed0
		x"034c197c", -- 7ed4
		x"00030343", -- 7ed8
		x"6100feec", -- 7edc
		x"660000ca", -- 7ee0
		x"2a2c035c", -- 7ee4
		x"41f8fdd2", -- 7ee8
		x"42305000", -- 7eec
		x"4a866730", -- 7ef0
		x"6d180c86", -- 7ef4
		x"00000002", -- 7ef8
		x"673c0c86", -- 7efc
		x"00000003", -- 7f00
		x"67343b7c", -- 7f04
		x"fffffff2", -- 7f08
		x"60164a10", -- 7f0c
		x"67084eba", -- 7f10
		x"023c41f8", -- 7f14
		x"fdd26100", -- 7f18
		x"00aa3b7c", -- 7f1c
		x"0001fff2", -- 7f20
		x"4a106704", -- 7f24
		x"610001a8", -- 7f28
		x"0c86ffff", -- 7f2c
		x"fffc6600", -- 7f30
		x"ff2e6000", -- 7f34
		x"00740c07", -- 7f38
		x"00016600", -- 7f3c
		x"006c4a10", -- 7f40
		x"67000066", -- 7f44
		x"61000188", -- 7f48
		x"41f8fdd2", -- 7f4c
		x"4ebad87a", -- 7f50
		x"007c0700", -- 7f54
		x"197c0001", -- 7f58
		x"00ba197c", -- 7f5c
		x"000000bb", -- 7f60
		x"08ac0000", -- 7f64
		x"00c008ac", -- 7f68
		x"000200c0", -- 7f6c
		x"08ec0002", -- 7f70
		x"000b08ac", -- 7f74
		x"0006000a", -- 7f78
		x"56e7027c", -- 7f7c
		x"f0ff082c", -- 7f80
		x"0002000b", -- 7f84
		x"66f84a1f", -- 7f88
		x"670608ec", -- 7f8c
		x"0006000a", -- 7f90
		x"41f8fdd2", -- 7f94
		x"2948034c", -- 7f98
		x"0c060002", -- 7f9c
		x"6700fec0", -- 7fa0
		x"43e9fffc", -- 7fa4
		x"6000feb8", -- 7fa8
		x"08380007", -- 7fac
		x"fdcc6600", -- 7fb0
		x"fd264eba", -- 7fb4
		x"d79441fa", -- 7fb8
		x"d9dc6100", -- 7fbc
		x"d80c6000", -- 7fc0
		x"fd1608f8", -- 7fc4
		x"0005fdcc", -- 7fc8
		x"0c410100", -- 7fcc
		x"6702613a", -- 7fd0
		x"4e7548e7", -- 7fd4
		x"80c02078", -- 7fd8
		x"fed443e8", -- 7fdc
		x"00dc2149", -- 7fe0
		x"000c08f8", -- 7fe4
		x"0007feda", -- 7fe8
		x"701f4219", -- 7fec
		x"51c8fffc", -- 7ff0
		x"4cdf0301", -- 7ff4
		x"4e7548e7", -- 7ff8
		x"f8c0183c", -- 7ffc
		x"00ff6010", -- 8000
		x"48e7f8c0", -- 8004
		x"183c0001", -- 8008
		x"600648e7", -- 800c
		x"f8c04204", -- 8010
		x"2878fed4", -- 8014
		x"41ec00dc", -- 8018
		x"42801001", -- 801c
		x"760880c3", -- 8020
		x"41f00000", -- 8024
		x"48407607", -- 8028
		x"96404a04", -- 802c
		x"6d066608", -- 8030
		x"07906006", -- 8034
		x"07106002", -- 8038
		x"07d04cdf", -- 803c
		x"031f4e75", -- 8040
		x"0c070002", -- 8044
		x"672a0838", -- 8048
		x"0007fdcc", -- 804c
		x"6622302c", -- 8050
		x"0046e248", -- 8054
		x"5e402f01", -- 8058
		x"222dfff4", -- 805c
		x"52415240", -- 8060
		x"4eac003c", -- 8064
		x"10186706", -- 8068
		x"4eac0036", -- 806c
		x"60f6221f", -- 8070
		x"4e750c07", -- 8074
		x"000267f8", -- 8078
		x"08380007", -- 807c
		x"fdcc66f0", -- 8080
		x"5248302c", -- 8084
		x"0046e248", -- 8088
		x"61cc48e7", -- 808c
		x"c080296d", -- 8090
		x"fff40350", -- 8094
		x"41f8fdd2", -- 8098
		x"2948034c", -- 809c
		x"197c0002", -- 80a0
		x"03436100", -- 80a4
		x"fd22661e", -- 80a8
		x"103c0020", -- 80ac
		x"4eac0036", -- 80b0
		x"222c035c", -- 80b4
		x"60061018", -- 80b8
		x"4eac0036", -- 80bc
		x"51c9fff8", -- 80c0
		x"4cdf0103", -- 80c4
		x"4e754cdf", -- 80c8
		x"01036000", -- 80cc
		x"fedc0c07", -- 80d0
		x"0002679c", -- 80d4
		x"08380007", -- 80d8
		x"fdcc6694", -- 80dc
		x"2f01222d", -- 80e0
		x"fff852ad", -- 80e4
		x"fff8302c", -- 80e8
		x"00565540", -- 80ec
		x"b06dfffa", -- 80f0
		x"6c0a202d", -- 80f4
		x"fffc5480", -- 80f8
		x"2b40fff8", -- 80fc
		x"302c0046", -- 8100
		x"e2486000", -- 8104
		x"ff580c07", -- 8108
		x"00026700", -- 810c
		x"ff6448e7", -- 8110
		x"e000202d", -- 8114
		x"fffc5480", -- 8118
		x"2b40fff8", -- 811c
		x"322c0056", -- 8120
		x"5541302c", -- 8124
		x"0046e248", -- 8128
		x"52404eac", -- 812c
		x"003c7020", -- 8130
		x"342c0046", -- 8134
		x"e24a4eac", -- 8138
		x"00365342", -- 813c
		x"6ef85341", -- 8140
		x"b26dfffa", -- 8144
		x"66dc4cdf", -- 8148
		x"00074e75", -- 814c
		x"08380007", -- 8150
		x"fdcc6600", -- 8154
		x"ff1c48e7", -- 8158
		x"c0887001", -- 815c
		x"322c032e", -- 8160
		x"4eac003c", -- 8164
		x"526c032e", -- 8168
		x"302c0056", -- 816c
		x"5540b06c", -- 8170
		x"032e6c06", -- 8174
		x"397c0001", -- 8178
		x"032e322c", -- 817c
		x"0046e249", -- 8180
		x"10186708", -- 8184
		x"4eac0036", -- 8188
		x"53416ef4", -- 818c
		x"4cdf1103", -- 8190
		x"4e756000", -- 8194
		x"46266000", -- 8198
		x"49c46000", -- 819c
		x"46b64ef9", -- 81a0
		x"000198d0", -- 81a4
		x"4ef83242", -- 81a8
		x"4ef8323e", -- 81ac
		x"4ef831a6", -- 81b0
		x"4ef834da", -- 81b4
		x"4ef830fe", -- 81b8
		x"4ef8361e", -- 81bc
		x"4ef835b8", -- 81c0
		x"4ef83372", -- 81c4
		x"4ef83398", -- 81c8
		x"205f225f", -- 81cc
		x"245f7800", -- 81d0
		x"181f7000", -- 81d4
		x"10196718", -- 81d8
		x"7c001c12", -- 81dc
		x"3e06de40", -- 81e0
		x"be446e0e", -- 81e4
		x"14c745f2", -- 81e8
		x"600014d9", -- 81ec
		x"53406efa", -- 81f0
		x"4ed03b7c", -- 81f4
		x"fff8fffe", -- 81f8
		x"4e4a205f", -- 81fc
		x"201f6e08", -- 8200
		x"dffc0000", -- 8204
		x"00144ed0", -- 8208
		x"221f6fe6", -- 820c
		x"225f7400", -- 8210
		x"14115242", -- 8214
		x"2c01dc80", -- 8218
		x"b4866dd6", -- 821c
		x"3c1f261f", -- 8220
		x"6fd02c03", -- 8224
		x"dc80245f", -- 8228
		x"7800181f", -- 822c
		x"7e003e04", -- 8230
		x"5287be86", -- 8234
		x"6dbc7e00", -- 8238
		x"1e125287", -- 823c
		x"be836db2", -- 8240
		x"be466c04", -- 8244
		x"53461486", -- 8248
		x"43f11800", -- 824c
		x"45f23800", -- 8250
		x"b5c96e08", -- 8254
		x"14d95380", -- 8258
		x"6efa4ed0", -- 825c
		x"43f10000", -- 8260
		x"45f20000", -- 8264
		x"15215380", -- 8268
		x"6efa4ed0", -- 826c
		x"00004e56", -- 8270
		x"0000302d", -- 8274
		x"fffe48c0", -- 8278
		x"2f00487a", -- 827c
		x"00184eba", -- 8280
		x"ff304a1f", -- 8284
		x"66000006", -- 8288
		x"4ebadfba", -- 828c
		x"422e0008", -- 8290
		x"4e5e4e75", -- 8294
		x"00027000", -- 8298
		x"00004e56", -- 829c
		x"0000558f", -- 82a0
		x"4eba2772", -- 82a4
		x"301f48c0", -- 82a8
		x"2f00487a", -- 82ac
		x"000e4eba", -- 82b0
		x"ff001d5f", -- 82b4
		x"00084e5e", -- 82b8
		x"4e750006", -- 82bc
		x"40800000", -- 82c0
		x"80000000", -- 82c4
		x"4e560000", -- 82c8
		x"558f4eba", -- 82cc
		x"2748301f", -- 82d0
		x"02400007", -- 82d4
		x"7207b240", -- 82d8
		x"57c00200", -- 82dc
		x"00011d40", -- 82e0
		x"00084e5e", -- 82e4
		x"4e750000", -- 82e8
		x"4e56fff8", -- 82ec
		x"1d7c0001", -- 82f0
		x"00142d79", -- 82f4
		x"fffffed4", -- 82f8
		x"fff84a2e", -- 82fc
		x"00126600", -- 8300
		x"0022206e", -- 8304
		x"fff8226e", -- 8308
		x"000c7000", -- 830c
		x"10280060", -- 8310
		x"3280226e", -- 8314
		x"00087000", -- 8318
		x"10280061", -- 831c
		x"32806000", -- 8320
		x"017a2f2d", -- 8324
		x"fff62f0e", -- 8328
		x"487a0160", -- 832c
		x"2b4ffff6", -- 8330
		x"206efff8", -- 8334
		x"0228ff1f", -- 8338
		x"005e7000", -- 833c
		x"eb888128", -- 8340
		x"005e0228", -- 8344
		x"00e0005e", -- 8348
		x"701f8128", -- 834c
		x"005e117c", -- 8350
		x"0000005f", -- 8354
		x"226e000c", -- 8358
		x"11690001", -- 835c
		x"0060226e", -- 8360
		x"00081169", -- 8364
		x"00010061", -- 8368
		x"558f4eba", -- 836c
		x"26a84a5f", -- 8370
		x"6600000a", -- 8374
		x"3b7c0001", -- 8378
		x"fffe4e4a", -- 837c
		x"558f4eba", -- 8380
		x"ff1a4a1f", -- 8384
		x"67000014", -- 8388
		x"4eba5364", -- 838c
		x"558f4eba", -- 8390
		x"53683d5f", -- 8394
		x"fffe6000", -- 8398
		x"0034558f", -- 839c
		x"4ebaff26", -- 83a0
		x"4a1f6700", -- 83a4
		x"0010558f", -- 83a8
		x"4eba538a", -- 83ac
		x"3d5ffffe", -- 83b0
		x"6000001a", -- 83b4
		x"206e0008", -- 83b8
		x"4a506700", -- 83bc
		x"000a3b7c", -- 83c0
		x"0001fffe", -- 83c4
		x"4e4a3d7c", -- 83c8
		x"fffffffe", -- 83cc
		x"3d7cffff", -- 83d0
		x"fffc526e", -- 83d4
		x"fffc206e", -- 83d8
		x"fff80228", -- 83dc
		x"ffe0005e", -- 83e0
		x"302efffc", -- 83e4
		x"8128005e", -- 83e8
		x"558f558f", -- 83ec
		x"4eba2626", -- 83f0
		x"3f2efffe", -- 83f4
		x"4eba516e", -- 83f8
		x"4a1f6700", -- 83fc
		x"00066000", -- 8400
		x"00220c6e", -- 8404
		x"001ffffc", -- 8408
		x"6dc8206e", -- 840c
		x"fff80228", -- 8410
		x"ffe0005e", -- 8414
		x"701f8128", -- 8418
		x"005e3b7c", -- 841c
		x"0001fffe", -- 8420
		x"4e4a558f", -- 8424
		x"206efff8", -- 8428
		x"48680072", -- 842c
		x"226e000c", -- 8430
		x"3f11226e", -- 8434
		x"00083f11", -- 8438
		x"4eba257e", -- 843c
		x"4a1f6600", -- 8440
		x"003c206e", -- 8444
		x"00084a50", -- 8448
		x"57c0122e", -- 844c
		x"00100841", -- 8450
		x"0000c001", -- 8454
		x"6700000a", -- 8458
		x"3b7c0001", -- 845c
		x"fffe4e4a", -- 8460
		x"4eba510c", -- 8464
		x"206efff8", -- 8468
		x"48680072", -- 846c
		x"226e000c", -- 8470
		x"3f11226e", -- 8474
		x"00083f11", -- 8478
		x"4eba2532", -- 847c
		x"2b6f0008", -- 8480
		x"fff6defc", -- 8484
		x"000c4efa", -- 8488
		x"00122c5f", -- 848c
		x"2b5ffff6", -- 8490
		x"558f4eba", -- 8494
		x"fdda1d5f", -- 8498
		x"00144e5e", -- 849c
		x"205fdefc", -- 84a0
		x"000c4ed0", -- 84a4
		x"00014e56", -- 84a8
		x"00002079", -- 84ac
		x"fffffed4", -- 84b0
		x"226e0008", -- 84b4
		x"24690010", -- 84b8
		x"24a8005e", -- 84bc
		x"558f4eba", -- 84c0
		x"fdda558f", -- 84c4
		x"4ebafdfe", -- 84c8
		x"101f801f", -- 84cc
		x"66000010", -- 84d0
		x"206e0008", -- 84d4
		x"22680010", -- 84d8
		x"137c00ff", -- 84dc
		x"0003206e", -- 84e0
		x"00082268", -- 84e4
		x"000c12bc", -- 84e8
		x"00014e5e", -- 84ec
		x"2e9f4e75", -- 84f0
		x"00004e56", -- 84f4
		x"fff8422e", -- 84f8
		x"00202d79", -- 84fc
		x"fffffed4", -- 8500
		x"fff8206e", -- 8504
		x"001c4a10", -- 8508
		x"66000034", -- 850c
		x"206e001c", -- 8510
		x"10bc0001", -- 8514
		x"206efff8", -- 8518
		x"1028005f", -- 851c
		x"02800000", -- 8520
		x"000f226e", -- 8524
		x"00183280", -- 8528
		x"1028005f", -- 852c
		x"e8880280", -- 8530
		x"0000000f", -- 8534
		x"226e0014", -- 8538
		x"32806000", -- 853c
		x"0170206e", -- 8540
		x"fff8226e", -- 8544
		x"00180228", -- 8548
		x"00f0005f", -- 854c
		x"30118128", -- 8550
		x"005f226e", -- 8554
		x"00140228", -- 8558
		x"000f005f", -- 855c
		x"3011e988", -- 8560
		x"8128005f", -- 8564
		x"70001028", -- 8568
		x"0060e940", -- 856c
		x"226e0018", -- 8570
		x"d0513d40", -- 8574
		x"fffe558f", -- 8578
		x"486800fc", -- 857c
		x"3f2efffe", -- 8580
		x"70001028", -- 8584
		x"00613f00", -- 8588
		x"4eba242e", -- 858c
		x"102e000a", -- 8590
		x"c01f6600", -- 8594
		x"01182f2d", -- 8598
		x"fff62f0e", -- 859c
		x"487a00b8", -- 85a0
		x"2b4ffff6", -- 85a4
		x"206efff8", -- 85a8
		x"0228ff1f", -- 85ac
		x"005e7000", -- 85b0
		x"eb888128", -- 85b4
		x"005e4eba", -- 85b8
		x"4fbc206e", -- 85bc
		x"000c4a10", -- 85c0
		x"66000008", -- 85c4
		x"2f0e4eba", -- 85c8
		x"fede4879", -- 85cc
		x"fffffdd2", -- 85d0
		x"2f3c0000", -- 85d4
		x"010042a7", -- 85d8
		x"4eba4fa2", -- 85dc
		x"206e0014", -- 85e0
		x"7007b050", -- 85e4
		x"57c0c02e", -- 85e8
		x"000a6700", -- 85ec
		x"001a206e", -- 85f0
		x"fff84868", -- 85f4
		x"00fc3f2e", -- 85f8
		x"fffe7000", -- 85fc
		x"10280061", -- 8600
		x"3f004eba", -- 8604
		x"23a83d7c", -- 8608
		x"fffffffc", -- 860c
		x"526efffc", -- 8610
		x"206efff8", -- 8614
		x"0228ff1f", -- 8618
		x"005e302e", -- 861c
		x"fffceb88", -- 8620
		x"8128005e", -- 8624
		x"558f4eba", -- 8628
		x"4eda4a1f", -- 862c
		x"67000012", -- 8630
		x"2f0e4eba", -- 8634
		x"fe721d7c", -- 8638
		x"fe010020", -- 863c
		x"6000000a", -- 8640
		x"0c6e0006", -- 8644
		x"fffc6dc4", -- 8648
		x"2b6f0008", -- 864c
		x"fff6defc", -- 8650
		x"000c4efa", -- 8654
		x"00582c5f", -- 8658
		x"2b5ffff6", -- 865c
		x"4a2e0008", -- 8660
		x"67000040", -- 8664
		x"7003b06d", -- 8668
		x"fffe6600", -- 866c
		x"000e206e", -- 8670
		x"001430bc", -- 8674
		x"00076000", -- 8678
		x"002a7001", -- 867c
		x"b06dfffe", -- 8680
		x"57c0c02e", -- 8684
		x"000a6700", -- 8688
		x"001a206e", -- 868c
		x"fff84868", -- 8690
		x"00fc3f2e", -- 8694
		x"fffe7000", -- 8698
		x"10280061", -- 869c
		x"3f004eba", -- 86a0
		x"230c558f", -- 86a4
		x"4ebafbc8", -- 86a8
		x"1d5f0020", -- 86ac
		x"4e5e205f", -- 86b0
		x"defc0018", -- 86b4
		x"4ed00000", -- 86b8
		x"4e56fff8", -- 86bc
		x"7001b06e", -- 86c0
		x"001e6700", -- 86c4
		x"000a422e", -- 86c8
		x"00206000", -- 86cc
		x"00a42079", -- 86d0
		x"fffffed4", -- 86d4
		x"41e8005e", -- 86d8
		x"2d48fff8", -- 86dc
		x"206e001a", -- 86e0
		x"4a106700", -- 86e4
		x"0024206e", -- 86e8
		x"fff80210", -- 86ec
		x"ffe0302e", -- 86f0
		x"00188110", -- 86f4
		x"226e0014", -- 86f8
		x"11690001", -- 86fc
		x"0002117c", -- 8700
		x"00000003", -- 8704
		x"60000012", -- 8708
		x"206efff8", -- 870c
		x"226e0014", -- 8710
		x"70001028", -- 8714
		x"00023280", -- 8718
		x"206e0010", -- 871c
		x"30100240", -- 8720
		x"000f3d40", -- 8724
		x"fffe206e", -- 8728
		x"00103010", -- 872c
		x"6c04d07c", -- 8730
		x"000fe840", -- 8734
		x"3d40fffc", -- 8738
		x"558f2f2e", -- 873c
		x"001a486e", -- 8740
		x"fffe486e", -- 8744
		x"fffc2f2e", -- 8748
		x"000c2f2e", -- 874c
		x"00084227", -- 8750
		x"42274eba", -- 8754
		x"fd9e1d5f", -- 8758
		x"0020302e", -- 875c
		x"fffc48c0", -- 8760
		x"e980322e", -- 8764
		x"fffe48c1", -- 8768
		x"d081206e", -- 876c
		x"00103080", -- 8770
		x"4e5e205f", -- 8774
		x"defc0018", -- 8778
		x"4ed00000", -- 877c
		x"4e56fff4", -- 8780
		x"7001b06e", -- 8784
		x"001457c0", -- 8788
		x"c02e0012", -- 878c
		x"6700005e", -- 8790
		x"3d7cffff", -- 8794
		x"fffc526e", -- 8798
		x"fffc2d79", -- 879c
		x"fffffed4", -- 87a0
		x"fff4206e", -- 87a4
		x"fff4302e", -- 87a8
		x"fffc4230", -- 87ac
		x"00724a2e", -- 87b0
		x"00086700", -- 87b4
		x"00303d7c", -- 87b8
		x"fffffff8", -- 87bc
		x"526efff8", -- 87c0
		x"206efff4", -- 87c4
		x"302efffc", -- 87c8
		x"48c0e980", -- 87cc
		x"322efff8", -- 87d0
		x"48c1d081", -- 87d4
		x"43e800fc", -- 87d8
		x"42310800", -- 87dc
		x"0c6e000f", -- 87e0
		x"fff86dd8", -- 87e4
		x"0c6e001f", -- 87e8
		x"fffc6daa", -- 87ec
		x"1d7c0001", -- 87f0
		x"00163d7c", -- 87f4
		x"fffffffc", -- 87f8
		x"526efffc", -- 87fc
		x"3d7cffff", -- 8800
		x"fffe526e", -- 8804
		x"fffe558f", -- 8808
		x"1f2e0012", -- 880c
		x"1f3c0001", -- 8810
		x"486efffc", -- 8814
		x"486efffe", -- 8818
		x"4ebaface", -- 881c
		x"4a1f6700", -- 8820
		x"004e3d7c", -- 8824
		x"fffffff8", -- 8828
		x"526efff8", -- 882c
		x"3d7cffff", -- 8830
		x"fffa526e", -- 8834
		x"fffa558f", -- 8838
		x"486e0012", -- 883c
		x"486efff8", -- 8840
		x"486efffa", -- 8844
		x"2f2e000e", -- 8848
		x"2f2e000a", -- 884c
		x"1f2e0008", -- 8850
		x"1f3c0001", -- 8854
		x"4ebafc9c", -- 8858
		x"4a1f6700", -- 885c
		x"00066000", -- 8860
		x"00224a6e", -- 8864
		x"fffa6dca", -- 8868
		x"4a6efff8", -- 886c
		x"6dba4a6e", -- 8870
		x"fffe6d8e", -- 8874
		x"701fb06e", -- 8878
		x"fffc6e00", -- 887c
		x"ff7c422e", -- 8880
		x"00164e5e", -- 8884
		x"205fdefc", -- 8888
		x"000e4ed0", -- 888c
		x"00004e56", -- 8890
		x"fff81d7c", -- 8894
		x"00010016", -- 8898
		x"3d7cffff", -- 889c
		x"fffc526e", -- 88a0
		x"fffc3d7c", -- 88a4
		x"fffffffe", -- 88a8
		x"526efffe", -- 88ac
		x"558f1f2e", -- 88b0
		x"00124227", -- 88b4
		x"486efffc", -- 88b8
		x"486efffe", -- 88bc
		x"4ebafa2a", -- 88c0
		x"4a1f6700", -- 88c4
		x"006c3d7c", -- 88c8
		x"fffffff8", -- 88cc
		x"526efff8", -- 88d0
		x"3d7cffff", -- 88d4
		x"fffa526e", -- 88d8
		x"fffa4a6e", -- 88dc
		x"fffe57c0", -- 88e0
		x"4a6efff8", -- 88e4
		x"57c1c200", -- 88e8
		x"4a6efffa", -- 88ec
		x"57c0c001", -- 88f0
		x"6600002e", -- 88f4
		x"558f486e", -- 88f8
		x"0012486e", -- 88fc
		x"fff8486e", -- 8900
		x"fffa2f2e", -- 8904
		x"000e2f2e", -- 8908
		x"000a1f2e", -- 890c
		x"00081f3c", -- 8910
		x"00014eba", -- 8914
		x"fbde4a1f", -- 8918
		x"67000006", -- 891c
		x"6000002a", -- 8920
		x"7007b06e", -- 8924
		x"fffa6eae", -- 8928
		x"700fb06e", -- 892c
		x"fff86e9c", -- 8930
		x"7007b06e", -- 8934
		x"fffe6e00", -- 8938
		x"ff70701f", -- 893c
		x"b06efffc", -- 8940
		x"6e00ff5c", -- 8944
		x"422e0016", -- 8948
		x"4e5e205f", -- 894c
		x"defc000e", -- 8950
		x"4ed00000", -- 8954
		x"4e56fffc", -- 8958
		x"426efffe", -- 895c
		x"3d7c00ff", -- 8960
		x"fffc558f", -- 8964
		x"3f2e0014", -- 8968
		x"486e0012", -- 896c
		x"4267486e", -- 8970
		x"fffc486e", -- 8974
		x"fffe2f2e", -- 8978
		x"000e2f2e", -- 897c
		x"000a4eba", -- 8980
		x"fd381d5f", -- 8984
		x"00164e5e", -- 8988
		x"205fdefc", -- 898c
		x"000e4ed0", -- 8990
		x"00004e56", -- 8994
		x"fffc1d7c", -- 8998
		x"00010016", -- 899c
		x"3d7c00ff", -- 89a0
		x"fffc426e", -- 89a4
		x"fffe526e", -- 89a8
		x"fffe558f", -- 89ac
		x"3f2e0014", -- 89b0
		x"486e0012", -- 89b4
		x"4267486e", -- 89b8
		x"fffc486e", -- 89bc
		x"fffe2f2e", -- 89c0
		x"000e2f2e", -- 89c4
		x"000a4eba", -- 89c8
		x"fcf04a1f", -- 89cc
		x"67000006", -- 89d0
		x"60000014", -- 89d4
		x"1039ffff", -- 89d8
		x"fed84880", -- 89dc
		x"b06efffe", -- 89e0
		x"6ec4422e", -- 89e4
		x"00164e5e", -- 89e8
		x"205fdefc", -- 89ec
		x"000e4ed0", -- 89f0
		x"00004e56", -- 89f4
		x"fffc426e", -- 89f8
		x"fffe3d7c", -- 89fc
		x"00fffffc", -- 8a00
		x"558f3f2e", -- 8a04
		x"0014486e", -- 8a08
		x"00123f3c", -- 8a0c
		x"0014486e", -- 8a10
		x"fffc486e", -- 8a14
		x"fffe2f2e", -- 8a18
		x"000e2f2e", -- 8a1c
		x"000a4eba", -- 8a20
		x"fc981d5f", -- 8a24
		x"00164e5e", -- 8a28
		x"205fdefc", -- 8a2c
		x"000e4ed0", -- 8a30
		x"00004e56", -- 8a34
		x"fffa1d7c", -- 8a38
		x"00010016", -- 8a3c
		x"3d7c00ff", -- 8a40
		x"fffa2079", -- 8a44
		x"fffffed4", -- 8a48
		x"70001028", -- 8a4c
		x"005f3d40", -- 8a50
		x"fffe426e", -- 8a54
		x"fffc526e", -- 8a58
		x"fffc558f", -- 8a5c
		x"3f2e0014", -- 8a60
		x"486e0012", -- 8a64
		x"3f3c0014", -- 8a68
		x"486efffa", -- 8a6c
		x"486efffc", -- 8a70
		x"2f2e000e", -- 8a74
		x"2f2e000a", -- 8a78
		x"4ebafc3e", -- 8a7c
		x"4a1f6700", -- 8a80
		x"00066000", -- 8a84
		x"001e302e", -- 8a88
		x"fffcb06e", -- 8a8c
		x"fffe6700", -- 8a90
		x"00066000", -- 8a94
		x"000a0c6e", -- 8a98
		x"00fffffc", -- 8a9c
		x"6db8422e", -- 8aa0
		x"00164e5e", -- 8aa4
		x"205fdefc", -- 8aa8
		x"000e4ed0", -- 8aac
		x"00004e56", -- 8ab0
		x"fffc3d7c", -- 8ab4
		x"001efffc", -- 8ab8
		x"3d7c00ff", -- 8abc
		x"fffe558f", -- 8ac0
		x"3f2e0014", -- 8ac4
		x"486e0012", -- 8ac8
		x"3f3c0016", -- 8acc
		x"486efffc", -- 8ad0
		x"486efffe", -- 8ad4
		x"2f2e000e", -- 8ad8
		x"2f2e000a", -- 8adc
		x"4ebafbda", -- 8ae0
		x"1d5f0016", -- 8ae4
		x"4e5e205f", -- 8ae8
		x"defc000e", -- 8aec
		x"4ed00000", -- 8af0
		x"4e56fffc", -- 8af4
		x"1d7c0001", -- 8af8
		x"00163d7c", -- 8afc
		x"00fffffe", -- 8b00
		x"3d7cffff", -- 8b04
		x"fffc526e", -- 8b08
		x"fffc701e", -- 8b0c
		x"b06efffc", -- 8b10
		x"6700002e", -- 8b14
		x"558f3f2e", -- 8b18
		x"0014486e", -- 8b1c
		x"00123f3c", -- 8b20
		x"0016486e", -- 8b24
		x"fffc486e", -- 8b28
		x"fffe2f2e", -- 8b2c
		x"000e2f2e", -- 8b30
		x"000a4eba", -- 8b34
		x"fb844a1f", -- 8b38
		x"67000006", -- 8b3c
		x"6000000e", -- 8b40
		x"701fb06e", -- 8b44
		x"fffc6ebe", -- 8b48
		x"422e0016", -- 8b4c
		x"4e5e205f", -- 8b50
		x"defc000e", -- 8b54
		x"4ed00000", -- 8b58
		x"4e56fff2", -- 8b5c
		x"2f2dfff6", -- 8b60
		x"2f0e487a", -- 8b64
		x"00382b4f", -- 8b68
		x"fff63d7c", -- 8b6c
		x"e942fffe", -- 8b70
		x"558f2f2e", -- 8b74
		x"0008486e", -- 8b78
		x"fffe486e", -- 8b7c
		x"fff6486e", -- 8b80
		x"fffa486e", -- 8b84
		x"fff24eba", -- 8b88
		x"497e1d5f", -- 8b8c
		x"000c2b6f", -- 8b90
		x"0008fff6", -- 8b94
		x"defc000c", -- 8b98
		x"4efa0010", -- 8b9c
		x"2c5f2b5f", -- 8ba0
		x"fff64eba", -- 8ba4
		x"d6a0422e", -- 8ba8
		x"000c4e5e", -- 8bac
		x"2e9f4e75", -- 8bb0
		x"4e75e108", -- 8bb4
		x"1500e108", -- 8bb8
		x"00000000", -- 8bbc
		x"4e560000", -- 8bc0
		x"206e000a", -- 8bc4
		x"302e0008", -- 8bc8
		x"2f1048c0", -- 8bcc
		x"d1977000", -- 8bd0
		x"205f1010", -- 8bd4
		x"3d40000e", -- 8bd8
		x"4e5e205f", -- 8bdc
		x"5c4f4ed0", -- 8be0
		x"00004e56", -- 8be4
		x"fff0422e", -- 8be8
		x"000e7020", -- 8bec
		x"b06e0008", -- 8bf0
		x"5ec02079", -- 8bf4
		x"fffffed4", -- 8bf8
		x"322e0008", -- 8bfc
		x"3401e842", -- 8c00
		x"e34a0241", -- 8c04
		x"000f41e8", -- 8c08
		x"00dc2630", -- 8c0c
		x"2000e3ab", -- 8c10
		x"721fe2ab", -- 8c14
		x"c0036700", -- 8c18
		x"01022d6e", -- 8c1c
		x"000afff4", -- 8c20
		x"2f3c0001", -- 8c24
		x"0000302e", -- 8c28
		x"00080240", -- 8c2c
		x"001f48c0", -- 8c30
		x"2f004eba", -- 8c34
		x"f5780697", -- 8c38
		x"00600000", -- 8c3c
		x"206efff4", -- 8c40
		x"209f42ae", -- 8c44
		x"fff852ae", -- 8c48
		x"fff8206e", -- 8c4c
		x"fff4202e", -- 8c50
		x"fff84230", -- 8c54
		x"08070cae", -- 8c58
		x"0000001a", -- 8c5c
		x"fff86de6", -- 8c60
		x"558f2f2e", -- 8c64
		x"000a3f3c", -- 8c68
		x"00014eba", -- 8c6c
		x"ff50301f", -- 8c70
		x"48c02d40", -- 8c74
		x"fff8202e", -- 8c78
		x"fff80280", -- 8c7c
		x"0000007f", -- 8c80
		x"2d40fff8", -- 8c84
		x"7034b0ae", -- 8c88
		x"fff86600", -- 8c8c
		x"008e558f", -- 8c90
		x"2f2e000a", -- 8c94
		x"3f3c4009", -- 8c98
		x"4ebaff22", -- 8c9c
		x"558f2f2e", -- 8ca0
		x"000a3f3c", -- 8ca4
		x"400b4eba", -- 8ca8
		x"ff14301f", -- 8cac
		x"48c0e180", -- 8cb0
		x"321f48c1", -- 8cb4
		x"d0812d40", -- 8cb8
		x"fffc0cae", -- 8cbc
		x"00008000", -- 8cc0
		x"fffc6c00", -- 8cc4
		x"0056558f", -- 8cc8
		x"2f2e000a", -- 8ccc
		x"202efffc", -- 8cd0
		x"e3805280", -- 8cd4
		x"3f004eba", -- 8cd8
		x"fee4301f", -- 8cdc
		x"48c02d40", -- 8ce0
		x"fffc202e", -- 8ce4
		x"fffc0280", -- 8ce8
		x"0000007f", -- 8cec
		x"7201b280", -- 8cf0
		x"57c0558f", -- 8cf4
		x"2f2e000a", -- 8cf8
		x"3f3c402f", -- 8cfc
		x"2d40fff0", -- 8d00
		x"4ebafeba", -- 8d04
		x"202efff0", -- 8d08
		x"7203b25f", -- 8d0c
		x"57c1c200", -- 8d10
		x"67000008", -- 8d14
		x"1d7c0001", -- 8d18
		x"000e4e5e", -- 8d1c
		x"205f5c4f", -- 8d20
		x"4ed00000", -- 8d24
		x"4e56fffa", -- 8d28
		x"302dfffe", -- 8d2c
		x"48c02d40", -- 8d30
		x"fffc2f2d", -- 8d34
		x"fff62f0e", -- 8d38
		x"487a003a", -- 8d3c
		x"2b4ffff6", -- 8d40
		x"558f2f3c", -- 8d44
		x"00010000", -- 8d48
		x"202e0008", -- 8d4c
		x"02800000", -- 8d50
		x"001f2f00", -- 8d54
		x"4ebaf456", -- 8d58
		x"06970060", -- 8d5c
		x"00004eba", -- 8d60
		x"17481d5f", -- 8d64
		x"fffb2b6f", -- 8d68
		x"0008fff6", -- 8d6c
		x"defc000c", -- 8d70
		x"4efa0008", -- 8d74
		x"2c5f2b5f", -- 8d78
		x"fff63b6e", -- 8d7c
		x"fffefffe", -- 8d80
		x"4e4a4e5e", -- 8d84
		x"2e9f4e75", -- 8d88
		x"00004e56", -- 8d8c
		x"fff42d79", -- 8d90
		x"fffffed4", -- 8d94
		x"fff4206e", -- 8d98
		x"fff47012", -- 8d9c
		x"d0a80010", -- 8da0
		x"2d40fffc", -- 8da4
		x"7034d0a8", -- 8da8
		x"00102d40", -- 8dac
		x"fff8558f", -- 8db0
		x"2f2efffc", -- 8db4
		x"3f2e001a", -- 8db8
		x"4ebafe28", -- 8dbc
		x"4a1f6700", -- 8dc0
		x"00902f2d", -- 8dc4
		x"fff62f0e", -- 8dc8
		x"487a0078", -- 8dcc
		x"2b4ffff6", -- 8dd0
		x"206efff8", -- 8dd4
		x"116e0017", -- 8dd8
		x"0007206e", -- 8ddc
		x"fff84228", -- 8de0
		x"0008206e", -- 8de4
		x"fff84228", -- 8de8
		x"0009206e", -- 8dec
		x"fff84228", -- 8df0
		x"000a206e", -- 8df4
		x"fff8117c", -- 8df8
		x"ff07000b", -- 8dfc
		x"2f2efffc", -- 8e00
		x"206efff8", -- 8e04
		x"48680007", -- 8e08
		x"202e0010", -- 8e0c
		x"5a802f00", -- 8e10
		x"4eba184c", -- 8e14
		x"4aae000c", -- 8e18
		x"6f000012", -- 8e1c
		x"2f2efffc", -- 8e20
		x"2f2e0008", -- 8e24
		x"2f2e000c", -- 8e28
		x"4eba1834", -- 8e2c
		x"2f2efffc", -- 8e30
		x"4eba1978", -- 8e34
		x"2b6f0008", -- 8e38
		x"fff6defc", -- 8e3c
		x"000c4efa", -- 8e40
		x"00102c5f", -- 8e44
		x"2b5ffff6", -- 8e48
		x"2f2e0018", -- 8e4c
		x"4ebafed6", -- 8e50
		x"4e5e205f", -- 8e54
		x"defc0014", -- 8e58
		x"4ed00000", -- 8e5c
		x"4e56ffe8", -- 8e60
		x"2d79ffff", -- 8e64
		x"fed4fff0", -- 8e68
		x"206efff0", -- 8e6c
		x"7012d0a8", -- 8e70
		x"00102d40", -- 8e74
		x"fff87034", -- 8e78
		x"d0a80010", -- 8e7c
		x"2d40fff4", -- 8e80
		x"558f2f2e", -- 8e84
		x"fff83f2e", -- 8e88
		x"000e4eba", -- 8e8c
		x"fd564a1f", -- 8e90
		x"6700013a", -- 8e94
		x"2d6efff4", -- 8e98
		x"ffec206e", -- 8e9c
		x"ffec2d48", -- 8ea0
		x"ffe82f2d", -- 8ea4
		x"fff62f0e", -- 8ea8
		x"487a00b0", -- 8eac
		x"2b4ffff6", -- 8eb0
		x"206effe8", -- 8eb4
		x"7000721c", -- 8eb8
		x"6f0610c0", -- 8ebc
		x"53816efa", -- 8ec0
		x"7003b0ae", -- 8ec4
		x"00086700", -- 8ec8
		x"00222d7c", -- 8ecc
		x"0000008b", -- 8ed0
		x"fffc2f2e", -- 8ed4
		x"fff8202e", -- 8ed8
		x"fff45080", -- 8edc
		x"2f00486e", -- 8ee0
		x"fffc4eba", -- 8ee4
		x"18086000", -- 8ee8
		x"00522d7c", -- 8eec
		x"00000028", -- 8ef0
		x"fffc2f2e", -- 8ef4
		x"fff8202e", -- 8ef8
		x"fff45080", -- 8efc
		x"2f00486e", -- 8f00
		x"fffc4eba", -- 8f04
		x"17e8206e", -- 8f08
		x"ffe870fd", -- 8f0c
		x"b0a80010", -- 8f10
		x"57c07224", -- 8f14
		x"b2a8000c", -- 8f18
		x"5dc1c200", -- 8f1c
		x"6700001c", -- 8f20
		x"226effec", -- 8f24
		x"2d69001c", -- 8f28
		x"fffc2f2e", -- 8f2c
		x"fff82f28", -- 8f30
		x"0014486e", -- 8f34
		x"fffc4eba", -- 8f38
		x"17b4202e", -- 8f3c
		x"00084480", -- 8f40
		x"206effe8", -- 8f44
		x"b0a80010", -- 8f48
		x"6600ff66", -- 8f4c
		x"2b6f0008", -- 8f50
		x"fff6defc", -- 8f54
		x"000c4efa", -- 8f58
		x"00102c5f", -- 8f5c
		x"2b5ffff6", -- 8f60
		x"2f2e000c", -- 8f64
		x"4ebafdbe", -- 8f68
		x"206effe8", -- 8f6c
		x"4aa80018", -- 8f70
		x"6700005a", -- 8f74
		x"20280018", -- 8f78
		x"90bc0000", -- 8f7c
		x"79182f00", -- 8f80
		x"487a0052", -- 8f84
		x"4ebaf22a", -- 8f88
		x"4a1f6700", -- 8f8c
		x"000e3b7c", -- 8f90
		x"0001fffe", -- 8f94
		x"4e4a6000", -- 8f98
		x"0034206e", -- 8f9c
		x"ffe82028", -- 8fa0
		x"001890bc", -- 8fa4
		x"00007918", -- 8fa8
		x"2f00487a", -- 8fac
		x"00304eba", -- 8fb0
		x"f2004a1f", -- 8fb4
		x"6700000e", -- 8fb8
		x"3b7c0004", -- 8fbc
		x"fffe4e4a", -- 8fc0
		x"6000000a", -- 8fc4
		x"3b7c0006", -- 8fc8
		x"fffe4e4a", -- 8fcc
		x"4e5e205f", -- 8fd0
		x"504f4ed0", -- 8fd4
		x"00060000", -- 8fd8
		x"28000808", -- 8fdc
		x"00060000", -- 8fe0
		x"03f3a005", -- 8fe4
		x"00004e56", -- 8fe8
		x"fffc2d6e", -- 8fec
		x"0010fffc", -- 8ff0
		x"206efffc", -- 8ff4
		x"216e000c", -- 8ff8
		x"000c216e", -- 8ffc
		x"00080010", -- 9000
		x"42a80014", -- 9004
		x"4e5e205f", -- 9008
		x"defc000c", -- 900c
		x"4ed00000", -- 9010
		x"4e56fff8", -- 9014
		x"2d6e000c", -- 9018
		x"fffc206e", -- 901c
		x"fffc4290", -- 9020
		x"4cba1e0f", -- 9024
		x"004c48a8", -- 9028
		x"1e0f0004", -- 902c
		x"4cba1e0f", -- 9030
		x"004048a8", -- 9034
		x"1e0f0014", -- 9038
		x"217c0000", -- 903c
		x"00010024", -- 9040
		x"43e80028", -- 9044
		x"2d49fff8", -- 9048
		x"226efff8", -- 904c
		x"22ae0008", -- 9050
		x"42a90004", -- 9054
		x"42a90008", -- 9058
		x"42a9000c", -- 905c
		x"4cba1e0f", -- 9060
		x"001048a8", -- 9064
		x"1e0f0038", -- 9068
		x"4e5e205f", -- 906c
		x"504f4ed0", -- 9070
		x"20202020", -- 9074
		x"20202020", -- 9078
		x"20202020", -- 907c
		x"20202020", -- 9080
		x"00004e56", -- 9084
		x"fffc2d6e", -- 9088
		x"000cfffc", -- 908c
		x"206efffc", -- 9090
		x"20ae0008", -- 9094
		x"42a80004", -- 9098
		x"42680008", -- 909c
		x"4268000a", -- 90a0
		x"4cba1e0f", -- 90a4
		x"001048a8", -- 90a8
		x"1e0f000c", -- 90ac
		x"4e5e205f", -- 90b0
		x"504f4ed0", -- 90b4
		x"20202020", -- 90b8
		x"20202020", -- 90bc
		x"20202020", -- 90c0
		x"20202020", -- 90c4
		x"00004e56", -- 90c8
		x"ffea206e", -- 90cc
		x"00104a10", -- 90d0
		x"57c00200", -- 90d4
		x"00011d40", -- 90d8
		x"ffff4a2e", -- 90dc
		x"ffff6600", -- 90e0
		x"00e0206e", -- 90e4
		x"0010226e", -- 90e8
		x"00107000", -- 90ec
		x"1011722f", -- 90f0
		x"b2300000", -- 90f4
		x"6600000c", -- 90f8
		x"1d7c0001", -- 90fc
		x"ffff6000", -- 9100
		x"00c0206e", -- 9104
		x"0010702f", -- 9108
		x"b0280001", -- 910c
		x"66000018", -- 9110
		x"206e000c", -- 9114
		x"20bc0000", -- 9118
		x"00012d7c", -- 911c
		x"00000002", -- 9120
		x"fffa6000", -- 9124
		x"0032206e", -- 9128
		x"00084cba", -- 912c
		x"1e0f02f0", -- 9130
		x"48901e0f", -- 9134
		x"206e0008", -- 9138
		x"4cba1e0f", -- 913c
		x"02f248a8", -- 9140
		x"1e0f0010", -- 9144
		x"206e000c", -- 9148
		x"20bc0000", -- 914c
		x"00022d7c", -- 9150
		x"00000001", -- 9154
		x"fffa1d7c", -- 9158
		x"0001fffe", -- 915c
		x"206e0008", -- 9160
		x"226e000c", -- 9164
		x"20112f00", -- 9168
		x"2f3c0000", -- 916c
		x"00242d48", -- 9170
		x"fff24eba", -- 9174
		x"f038206e", -- 9178
		x"fff2201f", -- 917c
		x"41f008dc", -- 9180
		x"4cba1e0f", -- 9184
		x"02aa4890", -- 9188
		x"1e0f206e", -- 918c
		x"0008226e", -- 9190
		x"000c2011", -- 9194
		x"2f002f3c", -- 9198
		x"00000024", -- 919c
		x"2d48fff2", -- 91a0
		x"4ebaf00a", -- 91a4
		x"206efff2", -- 91a8
		x"201f41f0", -- 91ac
		x"08ec4cba", -- 91b0
		x"1e0f027c", -- 91b4
		x"48901e0f", -- 91b8
		x"2d7c0000", -- 91bc
		x"0001fff6", -- 91c0
		x"206e0010", -- 91c4
		x"70001010", -- 91c8
		x"b0aefffa", -- 91cc
		x"5cc0122e", -- 91d0
		x"ffff0841", -- 91d4
		x"0000c200", -- 91d8
		x"6700022a", -- 91dc
		x"4a2efffe", -- 91e0
		x"670000f8", -- 91e4
		x"206e0010", -- 91e8
		x"202efffa", -- 91ec
		x"722fb230", -- 91f0
		x"08006600", -- 91f4
		x"0070206e", -- 91f8
		x"000c5290", -- 91fc
		x"206e0008", -- 9200
		x"226e000c", -- 9204
		x"20112f00", -- 9208
		x"2f3c0000", -- 920c
		x"00242d48", -- 9210
		x"fff24eba", -- 9214
		x"ef98206e", -- 9218
		x"fff2201f", -- 921c
		x"41f008dc", -- 9220
		x"4cba1e0f", -- 9224
		x"020a4890", -- 9228
		x"1e0f206e", -- 922c
		x"0008226e", -- 9230
		x"000c2011", -- 9234
		x"2f002f3c", -- 9238
		x"00000024", -- 923c
		x"2d48fff2", -- 9240
		x"4ebaef6a", -- 9244
		x"206efff2", -- 9248
		x"201f41f0", -- 924c
		x"08ec4cba", -- 9250
		x"1e0f01dc", -- 9254
		x"48901e0f", -- 9258
		x"2d7c0000", -- 925c
		x"0001fff6", -- 9260
		x"60000074", -- 9264
		x"206e0010", -- 9268
		x"202efffa", -- 926c
		x"723cb230", -- 9270
		x"08006600", -- 9274
		x"0012422e", -- 9278
		x"fffe2d7c", -- 927c
		x"00000001", -- 9280
		x"fff66000", -- 9284
		x"00527011", -- 9288
		x"b0aefff6", -- 928c
		x"6f000042", -- 9290
		x"206e0010", -- 9294
		x"202efffa", -- 9298
		x"226e0008", -- 929c
		x"246e000c", -- 92a0
		x"22122f01", -- 92a4
		x"2f3c0000", -- 92a8
		x"002448ee", -- 92ac
		x"0301ffea", -- 92b0
		x"4ebaeefa", -- 92b4
		x"4cee0301", -- 92b8
		x"ffea221f", -- 92bc
		x"242efff6", -- 92c0
		x"d48113b0", -- 92c4
		x"080028db", -- 92c8
		x"52aefff6", -- 92cc
		x"60000008", -- 92d0
		x"1d7c0001", -- 92d4
		x"ffff6000", -- 92d8
		x"0124206e", -- 92dc
		x"0010202e", -- 92e0
		x"fffa722f", -- 92e4
		x"b2300800", -- 92e8
		x"6600000c", -- 92ec
		x"1d7c0001", -- 92f0
		x"ffff6000", -- 92f4
		x"0108206e", -- 92f8
		x"0010202e", -- 92fc
		x"fffa723e", -- 9300
		x"b2300800", -- 9304
		x"660000a6", -- 9308
		x"52aefffa", -- 930c
		x"206e0010", -- 9310
		x"70001010", -- 9314
		x"b0aefffa", -- 9318
		x"6d00008e", -- 931c
		x"206e0010", -- 9320
		x"202efffa", -- 9324
		x"722fb230", -- 9328
		x"08006700", -- 932c
		x"000c1d7c", -- 9330
		x"0001ffff", -- 9334
		x"60000072", -- 9338
		x"1d7c0001", -- 933c
		x"fffe206e", -- 9340
		x"000c5290", -- 9344
		x"206e0008", -- 9348
		x"226e000c", -- 934c
		x"20112f00", -- 9350
		x"2f3c0000", -- 9354
		x"00242d48", -- 9358
		x"fff24eba", -- 935c
		x"ee50206e", -- 9360
		x"fff2201f", -- 9364
		x"41f008dc", -- 9368
		x"4cba1e0f", -- 936c
		x"00c24890", -- 9370
		x"1e0f206e", -- 9374
		x"0008226e", -- 9378
		x"000c2011", -- 937c
		x"2f002f3c", -- 9380
		x"00000024", -- 9384
		x"2d48fff2", -- 9388
		x"4ebaee22", -- 938c
		x"206efff2", -- 9390
		x"201f41f0", -- 9394
		x"08ec4cba", -- 9398
		x"1e0f0094", -- 939c
		x"48901e0f", -- 93a0
		x"2d7c0000", -- 93a4
		x"0001fff6", -- 93a8
		x"60000052", -- 93ac
		x"7011b0ae", -- 93b0
		x"fff66f00", -- 93b4
		x"0042206e", -- 93b8
		x"0010202e", -- 93bc
		x"fffa226e", -- 93c0
		x"0008246e", -- 93c4
		x"000c2212", -- 93c8
		x"2f012f3c", -- 93cc
		x"00000024", -- 93d0
		x"48ee0301", -- 93d4
		x"ffea4eba", -- 93d8
		x"edd44cee", -- 93dc
		x"0301ffea", -- 93e0
		x"221f242e", -- 93e4
		x"fff6d481", -- 93e8
		x"13b00800", -- 93ec
		x"28eb52ae", -- 93f0
		x"fff66000", -- 93f4
		x"00081d7c", -- 93f8
		x"0001ffff", -- 93fc
		x"52aefffa", -- 9400
		x"6000fdbe", -- 9404
		x"102effff", -- 9408
		x"08400000", -- 940c
		x"02000001", -- 9410
		x"1d400014", -- 9414
		x"4e5e205f", -- 9418
		x"defc000c", -- 941c
		x"4ed05359", -- 9420
		x"5354454d", -- 9424
		x"53202020", -- 9428
		x"20202020", -- 942c
		x"20202020", -- 9430
		x"20202020", -- 9434
		x"20202020", -- 9438
		x"20202020", -- 943c
		x"20200000", -- 9440
		x"4e56fff8", -- 9444
		x"2079ffff", -- 9448
		x"fed47034", -- 944c
		x"d0a80010", -- 9450
		x"2d40fff8", -- 9454
		x"2f3c0000", -- 9458
		x"00242f2e", -- 945c
		x"00144eba", -- 9460
		x"ed4c2d5f", -- 9464
		x"fffc206e", -- 9468
		x"fff84850", -- 946c
		x"203c0000", -- 9470
		x"0080d0ae", -- 9474
		x"fffc2f00", -- 9478
		x"2f3c0000", -- 947c
		x"00104eba", -- 9480
		x"fb66206e", -- 9484
		x"fff8217c", -- 9488
		x"00000001", -- 948c
		x"0018216e", -- 9490
		x"0008001c", -- 9494
		x"42a80020", -- 9498
		x"48680024", -- 949c
		x"2f2e000c", -- 94a0
		x"4ebafb6e", -- 94a4
		x"206efff8", -- 94a8
		x"42a80088", -- 94ac
		x"4868006c", -- 94b0
		x"2f2e0014", -- 94b4
		x"4ebafbcc", -- 94b8
		x"2f2e001c", -- 94bc
		x"2f2e0018", -- 94c0
		x"2f3c0000", -- 94c4
		x"00802f2e", -- 94c8
		x"fffc2f2e", -- 94cc
		x"00104eba", -- 94d0
		x"f8ba2f2e", -- 94d4
		x"001c2f3c", -- 94d8
		x"00000010", -- 94dc
		x"4ebaf97e", -- 94e0
		x"4e5e205f", -- 94e4
		x"defc0018", -- 94e8
		x"4ed00000", -- 94ec
		x"4e56fffc", -- 94f0
		x"2079ffff", -- 94f4
		x"fed47034", -- 94f8
		x"d0a80010", -- 94fc
		x"2d40fffc", -- 9500
		x"206efffc", -- 9504
		x"48502f3c", -- 9508
		x"00000010", -- 950c
		x"2f3c0000", -- 9510
		x"03e84eba", -- 9514
		x"fad2206e", -- 9518
		x"fffc42a8", -- 951c
		x"00182f2e", -- 9520
		x"000c2f2e", -- 9524
		x"00082f3c", -- 9528
		x"00000010", -- 952c
		x"42a742a7", -- 9530
		x"4ebaf858", -- 9534
		x"4e5e205f", -- 9538
		x"504f4ed0", -- 953c
		x"00004e56", -- 9540
		x"fff82079", -- 9544
		x"fffffed4", -- 9548
		x"7034d0a8", -- 954c
		x"00102d40", -- 9550
		x"fff82f3c", -- 9554
		x"00000024", -- 9558
		x"2f2e0010", -- 955c
		x"4ebaec4e", -- 9560
		x"2d5ffffc", -- 9564
		x"206efff8", -- 9568
		x"4850203c", -- 956c
		x"00000084", -- 9570
		x"d0aefffc", -- 9574
		x"2f002f3c", -- 9578
		x"0000000e", -- 957c
		x"4ebafa68", -- 9580
		x"206efff8", -- 9584
		x"48680018", -- 9588
		x"2f2e0008", -- 958c
		x"4ebafa82", -- 9590
		x"206efff8", -- 9594
		x"48680060", -- 9598
		x"2f2e0010", -- 959c
		x"4ebafae4", -- 95a0
		x"206efff8", -- 95a4
		x"42a8007c", -- 95a8
		x"42a80080", -- 95ac
		x"217c0000", -- 95b0
		x"00010084", -- 95b4
		x"42a80088", -- 95b8
		x"4268008c", -- 95bc
		x"4268008e", -- 95c0
		x"2f2e0018", -- 95c4
		x"2f2e0014", -- 95c8
		x"2f3c0000", -- 95cc
		x"00842f2e", -- 95d0
		x"fffc2f2e", -- 95d4
		x"000c4eba", -- 95d8
		x"f7b22f2e", -- 95dc
		x"00182f3c", -- 95e0
		x"0000000e", -- 95e4
		x"4ebaf876", -- 95e8
		x"4e5e205f", -- 95ec
		x"defc0014", -- 95f0
		x"4ed00000", -- 95f4
		x"4e56fff4", -- 95f8
		x"2d79ffff", -- 95fc
		x"fed4fff8", -- 9600
		x"206efff8", -- 9604
		x"7034d0a8", -- 9608
		x"00102d40", -- 960c
		x"fffc2d6e", -- 9610
		x"fffcfff4", -- 9614
		x"226efff4", -- 9618
		x"48512f3c", -- 961c
		x"00000028", -- 9620
		x"2f3c0000", -- 9624
		x"00034eba", -- 9628
		x"f9be206e", -- 962c
		x"fff4216e", -- 9630
		x"00080014", -- 9634
		x"217c0000", -- 9638
		x"00010018", -- 963c
		x"216e0018", -- 9640
		x"001c216e", -- 9644
		x"00140020", -- 9648
		x"42a80024", -- 964c
		x"42a80028", -- 9650
		x"216e0010", -- 9654
		x"002c216e", -- 9658
		x"000c0030", -- 965c
		x"2f2e0020", -- 9660
		x"2f2e001c", -- 9664
		x"2f3c0000", -- 9668
		x"002842a7", -- 966c
		x"42a74eba", -- 9670
		x"f71a4e5e", -- 9674
		x"205fdefc", -- 9678
		x"001c4ed0", -- 967c
		x"00004e56", -- 9680
		x"fffc2079", -- 9684
		x"fffffed4", -- 9688
		x"7034d0a8", -- 968c
		x"00102d40", -- 9690
		x"fffc206e", -- 9694
		x"fffc4850", -- 9698
		x"2f3c0000", -- 969c
		x"00542f3c", -- 96a0
		x"00000016", -- 96a4
		x"4ebaf940", -- 96a8
		x"206efffc", -- 96ac
		x"48680018", -- 96b0
		x"2f2e0008", -- 96b4
		x"4ebaf95a", -- 96b8
		x"2f2e0010", -- 96bc
		x"2f2e000c", -- 96c0
		x"2f3c0000", -- 96c4
		x"005442a7", -- 96c8
		x"42a74eba", -- 96cc
		x"f6be2f2e", -- 96d0
		x"00102f3c", -- 96d4
		x"00000016", -- 96d8
		x"4ebaf782", -- 96dc
		x"4e5e205f", -- 96e0
		x"defc000c", -- 96e4
		x"4ed00000", -- 96e8
		x"4e56ffec", -- 96ec
		x"2f2dfff6", -- 96f0
		x"2f0e487a", -- 96f4
		x"00f42b4f", -- 96f8
		x"fff62d79", -- 96fc
		x"fffffed4", -- 9700
		x"fff4206e", -- 9704
		x"fff47012", -- 9708
		x"d0a80010", -- 970c
		x"2d40fffc", -- 9710
		x"7034d0a8", -- 9714
		x"00102d40", -- 9718
		x"fff8422e", -- 971c
		x"0008226e", -- 9720
		x"fffc237c", -- 9724
		x"0000ea60", -- 9728
		x"000442a8", -- 972c
		x"006e42a8", -- 9730
		x"006a43e8", -- 9734
		x"005e2d49", -- 9738
		x"fff0558f", -- 973c
		x"2f2efffc", -- 9740
		x"226efff0", -- 9744
		x"70001029", -- 9748
		x"00023f00", -- 974c
		x"4ebaf494", -- 9750
		x"4a1f6700", -- 9754
		x"00862d6e", -- 9758
		x"fff8ffec", -- 975c
		x"558f2f3c", -- 9760
		x"00010000", -- 9764
		x"206efff0", -- 9768
		x"10280002", -- 976c
		x"0200001f", -- 9770
		x"72001200", -- 9774
		x"2f014eba", -- 9778
		x"ea340697", -- 977c
		x"00600000", -- 9780
		x"4eba0d26", -- 9784
		x"4a1f6700", -- 9788
		x"0052206e", -- 978c
		x"fff07000", -- 9790
		x"10280002", -- 9794
		x"2f007000", -- 9798
		x"10280003", -- 979c
		x"2f004eba", -- 97a0
		x"fd4c206e", -- 97a4
		x"fff07000", -- 97a8
		x"10280002", -- 97ac
		x"2f007000", -- 97b0
		x"10280003", -- 97b4
		x"2f007000", -- 97b8
		x"10280001", -- 97bc
		x"2f004eba", -- 97c0
		x"febe206e", -- 97c4
		x"ffec4aa8", -- 97c8
		x"001857c0", -- 97cc
		x"c028001f", -- 97d0
		x"67000008", -- 97d4
		x"1d7c0001", -- 97d8
		x"00082b6f", -- 97dc
		x"0008fff6", -- 97e0
		x"defc000c", -- 97e4
		x"4efa0020", -- 97e8
		x"2c5f2b5f", -- 97ec
		x"fff6302d", -- 97f0
		x"fffe48c0", -- 97f4
		x"2f00487a", -- 97f8
		x"00124eba", -- 97fc
		x"e9b44a1f", -- 9800
		x"66000004", -- 9804
		x"4e4a4e5e", -- 9808
		x"4e750002", -- 980c
		x"60000001", -- 9810
		x"4e56fff4", -- 9814
		x"2d79ffff", -- 9818
		x"fed4fffc", -- 981c
		x"206efffc", -- 9820
		x"43e8005e", -- 9824
		x"2d49fff8", -- 9828
		x"226efff8", -- 982c
		x"70001029", -- 9830
		x"00022f00", -- 9834
		x"70001029", -- 9838
		x"00032f00", -- 983c
		x"246e0008", -- 9840
		x"2f2afff8", -- 9844
		x"2f2affdc", -- 9848
		x"70001029", -- 984c
		x"00012f00", -- 9850
		x"4ebafcec", -- 9854
		x"206e0008", -- 9858
		x"2d68ffe0", -- 985c
		x"fff42268", -- 9860
		x"000870ff", -- 9864
		x"b05157c0", -- 9868
		x"226efff4", -- 986c
		x"24680008", -- 9870
		x"3212b269", -- 9874
		x"002e57c1", -- 9878
		x"82006700", -- 987c
		x"0030246e", -- 9880
		x"fffc2569", -- 9884
		x"001c006e", -- 9888
		x"117c0001", -- 988c
		x"0018117c", -- 9890
		x"0001ffff", -- 9894
		x"26680010", -- 9898
		x"26a9003c", -- 989c
		x"2668000c", -- 98a0
		x"26a90030", -- 98a4
		x"26680008", -- 98a8
		x"36a9002e", -- 98ac
		x"4e5e2e9f", -- 98b0
		x"4e750000", -- 98b4
		x"4e56ffbc", -- 98b8
		x"422e0018", -- 98bc
		x"4eba04ae", -- 98c0
		x"422effff", -- 98c4
		x"2d79ffff", -- 98c8
		x"fed4ffd8", -- 98cc
		x"206effd8", -- 98d0
		x"43e8005e", -- 98d4
		x"2d49ffd4", -- 98d8
		x"7034d0a8", -- 98dc
		x"00102d40", -- 98e0
		x"ffe02d7c", -- 98e4
		x"fffffdd2", -- 98e8
		x"ffdc558f", -- 98ec
		x"2f2e0014", -- 98f0
		x"486efff8", -- 98f4
		x"2f2effdc", -- 98f8
		x"4ebaf7cc", -- 98fc
		x"4a1f6700", -- 9900
		x"02d4598f", -- 9904
		x"487a02d8", -- 9908
		x"2f2e0014", -- 990c
		x"4ebae8aa", -- 9910
		x"4a9f6600", -- 9914
		x"003a2f2d", -- 9918
		x"fff62f0e", -- 991c
		x"487a001a", -- 9920
		x"2b4ffff6", -- 9924
		x"2f0e4eba", -- 9928
		x"fee82b6f", -- 992c
		x"0008fff6", -- 9930
		x"defc000c", -- 9934
		x"4efa0014", -- 9938
		x"2c5f2b5f", -- 993c
		x"fff67004", -- 9940
		x"b06dfffe", -- 9944
		x"67000004", -- 9948
		x"4e4a6000", -- 994c
		x"0288206e", -- 9950
		x"ffd852a8", -- 9954
		x"006a2f2d", -- 9958
		x"fff62f0e", -- 995c
		x"487a0252", -- 9960
		x"2b4ffff6", -- 9964
		x"226effd4", -- 9968
		x"70001029", -- 996c
		x"00022f00", -- 9970
		x"70001029", -- 9974
		x"00032f00", -- 9978
		x"202efff8", -- 997c
		x"53802f00", -- 9980
		x"2f2effdc", -- 9984
		x"70001029", -- 9988
		x"00012f00", -- 998c
		x"2f28006a", -- 9990
		x"4ebafaae", -- 9994
		x"2d6effe0", -- 9998
		x"ffd0206e", -- 999c
		x"ffd043e8", -- 99a0
		x"00242d49", -- 99a4
		x"ffcc7001", -- 99a8
		x"b0a80020", -- 99ac
		x"6f00000c", -- 99b0
		x"1d7c0001", -- 99b4
		x"ffff6000", -- 99b8
		x"01ea206e", -- 99bc
		x"000870ff", -- 99c0
		x"b05057c0", -- 99c4
		x"206effcc", -- 99c8
		x"226e0008", -- 99cc
		x"3211b268", -- 99d0
		x"001a57c1", -- 99d4
		x"82006700", -- 99d8
		x"01ca1d7c", -- 99dc
		x"0001fffe", -- 99e0
		x"422efffd", -- 99e4
		x"426efff6", -- 99e8
		x"526efff6", -- 99ec
		x"4a2efffd", -- 99f0
		x"6600007c", -- 99f4
		x"206effdc", -- 99f8
		x"202efff8", -- 99fc
		x"2f002f3c", -- 9a00
		x"00000024", -- 9a04
		x"2d48ffc8", -- 9a08
		x"4ebae7a2", -- 9a0c
		x"206effc8", -- 9a10
		x"201f322e", -- 9a14
		x"fff648c1", -- 9a18
		x"d2804a30", -- 9a1c
		x"18db6600", -- 9a20
		x"000c1d7c", -- 9a24
		x"0001fffd", -- 9a28
		x"60000044", -- 9a2c
		x"206effcc", -- 9a30
		x"302efff6", -- 9a34
		x"226effdc", -- 9a38
		x"222efff8", -- 9a3c
		x"2f012f3c", -- 9a40
		x"00000024", -- 9a44
		x"48ee0301", -- 9a48
		x"ffbc4eba", -- 9a4c
		x"e7604cee", -- 9a50
		x"0301ffbc", -- 9a54
		x"221f342e", -- 9a58
		x"fff648c2", -- 9a5c
		x"d4811231", -- 9a60
		x"28dbb230", -- 9a64
		x"00ff6700", -- 9a68
		x"0006422e", -- 9a6c
		x"fffe0c6e", -- 9a70
		x"0010fff6", -- 9a74
		x"6d00ff72", -- 9a78
		x"4a2efffe", -- 9a7c
		x"67000124", -- 9a80
		x"206effdc", -- 9a84
		x"202efff8", -- 9a88
		x"2f002f3c", -- 9a8c
		x"00000024", -- 9a90
		x"2d48ffc8", -- 9a94
		x"4ebae716", -- 9a98
		x"206effc8", -- 9a9c
		x"201f41f0", -- 9aa0
		x"08dc4c90", -- 9aa4
		x"1e0f48ae", -- 9aa8
		x"1e0fffe4", -- 9aac
		x"206effcc", -- 9ab0
		x"226effdc", -- 9ab4
		x"202efff8", -- 9ab8
		x"2f002f3c", -- 9abc
		x"00000024", -- 9ac0
		x"48ee0300", -- 9ac4
		x"ffc44eba", -- 9ac8
		x"e6e44cee", -- 9acc
		x"0300ffc4", -- 9ad0
		x"201f43f1", -- 9ad4
		x"08dc4c90", -- 9ad8
		x"1c1f4891", -- 9adc
		x"1c1f7000", -- 9ae0
		x"226e0014", -- 9ae4
		x"10113d40", -- 9ae8
		x"fff6536e", -- 9aec
		x"fff6206e", -- 9af0
		x"0014302e", -- 9af4
		x"fff6722f", -- 9af8
		x"b2300000", -- 9afc
		x"57c04a6e", -- 9b00
		x"fff657c1", -- 9b04
		x"820067e2", -- 9b08
		x"7010d06e", -- 9b0c
		x"fff6206e", -- 9b10
		x"00141080", -- 9b14
		x"426efff4", -- 9b18
		x"526efff4", -- 9b1c
		x"206effcc", -- 9b20
		x"302efff4", -- 9b24
		x"226e0014", -- 9b28
		x"322efff6", -- 9b2c
		x"d26efff4", -- 9b30
		x"13b000ff", -- 9b34
		x"10000c6e", -- 9b38
		x"0010fff4", -- 9b3c
		x"6dda2f2d", -- 9b40
		x"fff62f0e", -- 9b44
		x"487a001a", -- 9b48
		x"2b4ffff6", -- 9b4c
		x"2f0e4eba", -- 9b50
		x"fcc02b6f", -- 9b54
		x"0008fff6", -- 9b58
		x"defc000c", -- 9b5c
		x"4efa0044", -- 9b60
		x"2c5f2b5f", -- 9b64
		x"fff67004", -- 9b68
		x"b06dfffe", -- 9b6c
		x"67000008", -- 9b70
		x"4e4a6000", -- 9b74
		x"002e206e", -- 9b78
		x"ffdc202e", -- 9b7c
		x"fff82f00", -- 9b80
		x"2f3c0000", -- 9b84
		x"00242d48", -- 9b88
		x"ffc84eba", -- 9b8c
		x"e620206e", -- 9b90
		x"ffc8201f", -- 9b94
		x"41f008dc", -- 9b98
		x"4cae1e0f", -- 9b9c
		x"ffe44890", -- 9ba0
		x"1e0f2b6f", -- 9ba4
		x"0008fff6", -- 9ba8
		x"defc000c", -- 9bac
		x"4efa001e", -- 9bb0
		x"2c5f2b5f", -- 9bb4
		x"fff67004", -- 9bb8
		x"b06dfffe", -- 9bbc
		x"6600000c", -- 9bc0
		x"1d7c0001", -- 9bc4
		x"ffff6000", -- 9bc8
		x"00044e4a", -- 9bcc
		x"4a2effff", -- 9bd0
		x"6700fd7c", -- 9bd4
		x"4e5e205f", -- 9bd8
		x"defc0010", -- 9bdc
		x"4ed00100", -- 9be0
		x"00004e56", -- 9be4
		x"ffe42d79", -- 9be8
		x"fffffed4", -- 9bec
		x"ffec206e", -- 9bf0
		x"ffec7034", -- 9bf4
		x"d0a80010", -- 9bf8
		x"2d40fff0", -- 9bfc
		x"4aa8006e", -- 9c00
		x"56c0122e", -- 9c04
		x"00080841", -- 9c08
		x"0000c001", -- 9c0c
		x"67000152", -- 9c10
		x"43e8005e", -- 9c14
		x"2d49ffe8", -- 9c18
		x"2d6efff0", -- 9c1c
		x"ffe442ae", -- 9c20
		x"fffc42ae", -- 9c24
		x"fff8202e", -- 9c28
		x"0012e180", -- 9c2c
		x"2d40fff4", -- 9c30
		x"0cae0000", -- 9c34
		x"0200000e", -- 9c38
		x"6f0000b8", -- 9c3c
		x"226effe8", -- 9c40
		x"70001029", -- 9c44
		x"00022f00", -- 9c48
		x"70001029", -- 9c4c
		x"00032f00", -- 9c50
		x"2f28006e", -- 9c54
		x"2f2efff8", -- 9c58
		x"2f3c0000", -- 9c5c
		x"02002f2e", -- 9c60
		x"fff42f2e", -- 9c64
		x"000a4eba", -- 9c68
		x"f98c2d7c", -- 9c6c
		x"00000200", -- 9c70
		x"fffc06ae", -- 9c74
		x"00000200", -- 9c78
		x"000a2d7c", -- 9c7c
		x"00000001", -- 9c80
		x"fff842ae", -- 9c84
		x"fff4202e", -- 9c88
		x"000e90ae", -- 9c8c
		x"fffc0c80", -- 9c90
		x"00000200", -- 9c94
		x"6f00005c", -- 9c98
		x"206effe8", -- 9c9c
		x"70001028", -- 9ca0
		x"00022f00", -- 9ca4
		x"70001028", -- 9ca8
		x"00032f00", -- 9cac
		x"226effec", -- 9cb0
		x"2f29006e", -- 9cb4
		x"2f2efff8", -- 9cb8
		x"2f3c0000", -- 9cbc
		x"02002f2e", -- 9cc0
		x"fff42f2e", -- 9cc4
		x"000a4eba", -- 9cc8
		x"f92c06ae", -- 9ccc
		x"00000200", -- 9cd0
		x"fffc06ae", -- 9cd4
		x"00000200", -- 9cd8
		x"000a206e", -- 9cdc
		x"ffe87000", -- 9ce0
		x"10280002", -- 9ce4
		x"2f002f3c", -- 9ce8
		x"00000003", -- 9cec
		x"4ebaf16e", -- 9cf0
		x"6094206e", -- 9cf4
		x"ffe87000", -- 9cf8
		x"10280002", -- 9cfc
		x"2f007000", -- 9d00
		x"10280003", -- 9d04
		x"2f00226e", -- 9d08
		x"ffec2f29", -- 9d0c
		x"006e2f2e", -- 9d10
		x"fff8202e", -- 9d14
		x"000e90ae", -- 9d18
		x"fffc2f00", -- 9d1c
		x"2f2efff4", -- 9d20
		x"2f2e000a", -- 9d24
		x"4ebaf8ce", -- 9d28
		x"206effe8", -- 9d2c
		x"70001028", -- 9d30
		x"00022f00", -- 9d34
		x"2f3c0000", -- 9d38
		x"00034eba", -- 9d3c
		x"f1200cae", -- 9d40
		x"00000200", -- 9d44
		x"000e6f00", -- 9d48
		x"0018206e", -- 9d4c
		x"ffe87000", -- 9d50
		x"10280002", -- 9d54
		x"2f002f3c", -- 9d58
		x"00000003", -- 9d5c
		x"4ebaf0fe", -- 9d60
		x"4e5e205f", -- 9d64
		x"defc000e", -- 9d68
		x"4ed00000", -- 9d6c
		x"4e56fffc", -- 9d70
		x"2079ffff", -- 9d74
		x"fed441e8", -- 9d78
		x"005e2d48", -- 9d7c
		x"fffc206e", -- 9d80
		x"fffc7000", -- 9d84
		x"10280002", -- 9d88
		x"2f007000", -- 9d8c
		x"10280003", -- 9d90
		x"2f004eba", -- 9d94
		x"f7584e5e", -- 9d98
		x"4e750000", -- 9d9c
		x"4e56ffe6", -- 9da0
		x"2f2dfff6", -- 9da4
		x"2f0e487a", -- 9da8
		x"01b22b4f", -- 9dac
		x"fff62d79", -- 9db0
		x"fffffed4", -- 9db4
		x"fff2206e", -- 9db8
		x"fff243e8", -- 9dbc
		x"005e2d49", -- 9dc0
		x"ffee7012", -- 9dc4
		x"d0a80010", -- 9dc8
		x"2d40fffa", -- 9dcc
		x"7034d0a8", -- 9dd0
		x"00102d40", -- 9dd4
		x"fff6226e", -- 9dd8
		x"000a4211", -- 9ddc
		x"4a2e0012", -- 9de0
		x"67000020", -- 9de4
		x"217aedcc", -- 9de8
		x"005e7001", -- 9dec
		x"b06e0014", -- 9df0
		x"57c0c02e", -- 9df4
		x"00086700", -- 9df8
		x"000642a8", -- 9dfc
		x"02fc6000", -- 9e00
		x"000c206e", -- 9e04
		x"fff2217a", -- 9e08
		x"edae005e", -- 9e0c
		x"558f2f2e", -- 9e10
		x"fffa206e", -- 9e14
		x"ffee7000", -- 9e18
		x"10280002", -- 9e1c
		x"3f004eba", -- 9e20
		x"edc24a1f", -- 9e24
		x"6700011e", -- 9e28
		x"1d7c0001", -- 9e2c
		x"ffff4a2e", -- 9e30
		x"00086700", -- 9e34
		x"0032206e", -- 9e38
		x"fff2226e", -- 9e3c
		x"ffee7000", -- 9e40
		x"10290002", -- 9e44
		x"3200e841", -- 9e48
		x"e3490240", -- 9e4c
		x"000f45e8", -- 9e50
		x"02fc2432", -- 9e54
		x"1000e1aa", -- 9e58
		x"701fe0aa", -- 9e5c
		x"4a826700", -- 9e60
		x"0006422e", -- 9e64
		x"ffff4a2e", -- 9e68
		x"ffff6700", -- 9e6c
		x"00d8206e", -- 9e70
		x"fff22028", -- 9e74
		x"005eb0ba", -- 9e78
		x"ed3a6600", -- 9e7c
		x"00c82d6e", -- 9e80
		x"fff6ffea", -- 9e84
		x"226effea", -- 9e88
		x"2d49ffe6", -- 9e8c
		x"246efffa", -- 9e90
		x"257c0000", -- 9e94
		x"13880004", -- 9e98
		x"246effee", -- 9e9c
		x"7000102a", -- 9ea0
		x"00022f00", -- 9ea4
		x"7000102a", -- 9ea8
		x"00032f00", -- 9eac
		x"4ebaf63e", -- 9eb0
		x"206effee", -- 9eb4
		x"70001028", -- 9eb8
		x"00022f00", -- 9ebc
		x"70001028", -- 9ec0
		x"00032f00", -- 9ec4
		x"70001028", -- 9ec8
		x"00012f00", -- 9ecc
		x"4ebaf7b0", -- 9ed0
		x"206effe6", -- 9ed4
		x"4aa80018", -- 9ed8
		x"57c0226e", -- 9edc
		x"ffeac029", -- 9ee0
		x"001f6700", -- 9ee4
		x"0060246e", -- 9ee8
		x"fff2266e", -- 9eec
		x"000e26aa", -- 9ef0
		x"005e558f", -- 9ef4
		x"4ebaf7f2", -- 9ef8
		x"206e000a", -- 9efc
		x"109f206e", -- 9f00
		x"000a102e", -- 9f04
		x"0008c010", -- 9f08
		x"6700003a", -- 9f0c
		x"206efff2", -- 9f10
		x"226effee", -- 9f14
		x"70001029", -- 9f18
		x"00023200", -- 9f1c
		x"e841e349", -- 9f20
		x"0240000f", -- 9f24
		x"45e802fc", -- 9f28
		x"74014400", -- 9f2c
		x"d03c021f", -- 9f30
		x"e1aa4682", -- 9f34
		x"c5b21000", -- 9f38
		x"74017600", -- 9f3c
		x"1602e1ab", -- 9f40
		x"87b21000", -- 9f44
		x"206e000a", -- 9f48
		x"1d500016", -- 9f4c
		x"2b6f0008", -- 9f50
		x"fff6defc", -- 9f54
		x"000c4efa", -- 9f58
		x"00262c5f", -- 9f5c
		x"2b5ffff6", -- 9f60
		x"422e0016", -- 9f64
		x"302dfffe", -- 9f68
		x"48c02f00", -- 9f6c
		x"487a001a", -- 9f70
		x"4ebae23e", -- 9f74
		x"4a1f6600", -- 9f78
		x"00064eba", -- 9f7c
		x"c2c84e5e", -- 9f80
		x"205fdefc", -- 9f84
		x"000e4ed0", -- 9f88
		x"00026000", -- 9f8c
		x"00004e56", -- 9f90
		x"ffea2f2d", -- 9f94
		x"fff62f0e", -- 9f98
		x"487a0414", -- 9f9c
		x"2b4ffff6", -- 9fa0
		x"2d79ffff", -- 9fa4
		x"fed4fff2", -- 9fa8
		x"206efff2", -- 9fac
		x"43e8005e", -- 9fb0
		x"2d49ffee", -- 9fb4
		x"7012d0a8", -- 9fb8
		x"00102d40", -- 9fbc
		x"fffa7034", -- 9fc0
		x"d0a80010", -- 9fc4
		x"2d40fff6", -- 9fc8
		x"226e000a", -- 9fcc
		x"42114a2e", -- 9fd0
		x"00126700", -- 9fd4
		x"0022217a", -- 9fd8
		x"ebde005e", -- 9fdc
		x"08a80003", -- 9fe0
		x"005c7001", -- 9fe4
		x"b06e0014", -- 9fe8
		x"57c0c02e", -- 9fec
		x"00086700", -- 9ff0
		x"000642a8", -- 9ff4
		x"02fc206e", -- 9ff8
		x"ffee7020", -- 9ffc
		x"b0280002", -- a000
		x"52c0226e", -- a004
		x"000a1211", -- a008
		x"08410000", -- a00c
		x"c2006700", -- a010
		x"03884a2e", -- a014
		x"00126700", -- a018
		x"000a422e", -- a01c
		x"00126000", -- a020
		x"0042206e", -- a024
		x"fff20828", -- a028
		x"0003005c", -- a02c
		x"56c04400", -- a030
		x"226effee", -- a034
		x"72001229", -- a038
		x"00033401", -- a03c
		x"e842e34a", -- a040
		x"0241000f", -- a044
		x"45e80092", -- a048
		x"26322000", -- a04c
		x"e3ab721f", -- a050
		x"e2ab0843", -- a054
		x"0000c600", -- a058
		x"67000008", -- a05c
		x"137c0018", -- a060
		x"0001206e", -- a064
		x"ffee7018", -- a068
		x"b0280001", -- a06c
		x"63000042", -- a070
		x"7008b028", -- a074
		x"00016600", -- a078
		x"000c117c", -- a07c
		x"00070001", -- a080
		x"6000002a", -- a084
		x"206effee", -- a088
		x"7007b028", -- a08c
		x"00016600", -- a090
		x"000c117c", -- a094
		x"00090001", -- a098
		x"60000012", -- a09c
		x"206effee", -- a0a0
		x"70001028", -- a0a4
		x"00015240", -- a0a8
		x"11400001", -- a0ac
		x"6000011c", -- a0b0
		x"206effee", -- a0b4
		x"117cff08", -- a0b8
		x"00017040", -- a0bc
		x"b0280003", -- a0c0
		x"63000050", -- a0c4
		x"206effee", -- a0c8
		x"70001028", -- a0cc
		x"00035240", -- a0d0
		x"11400003", -- a0d4
		x"226efff2", -- a0d8
		x"08290003", -- a0dc
		x"005c56c0", -- a0e0
		x"44000840", -- a0e4
		x"00007200", -- a0e8
		x"12280003", -- a0ec
		x"3401e842", -- a0f0
		x"e34a0241", -- a0f4
		x"000f45e9", -- a0f8
		x"00922632", -- a0fc
		x"2000e3ab", -- a100
		x"721fe2ab", -- a104
		x"8600703f", -- a108
		x"b0280003", -- a10c
		x"55c08003", -- a110
		x"67b2206e", -- a114
		x"ffee703f", -- a118
		x"b0280003", -- a11c
		x"640000ac", -- a120
		x"226efff2", -- a124
		x"08290003", -- a128
		x"005c56c0", -- a12c
		x"44004a00", -- a130
		x"67000048", -- a134
		x"4aa90092", -- a138
		x"56c04aa9", -- a13c
		x"009656c1", -- a140
		x"8200c22e", -- a144
		x"00086700", -- a148
		x"00327000", -- a14c
		x"10280002", -- a150
		x"3200e841", -- a154
		x"e3490240", -- a158
		x"000f45e9", -- a15c
		x"02fc7401", -- a160
		x"4400d03c", -- a164
		x"021fe1aa", -- a168
		x"4682c5b2", -- a16c
		x"10007401", -- a170
		x"76001602", -- a174
		x"e1ab87b2", -- a178
		x"1000206e", -- a17c
		x"fff208a8", -- a180
		x"0003005c", -- a184
		x"226effee", -- a188
		x"137cff00", -- a18c
		x"0003137c", -- a190
		x"ff080001", -- a194
		x"206effee", -- a198
		x"70001028", -- a19c
		x"00025240", -- a1a0
		x"11400002", -- a1a4
		x"701fb028", -- a1a8
		x"000255c0", -- a1ac
		x"558f2f2e", -- a1b0
		x"fffa7200", -- a1b4
		x"12280002", -- a1b8
		x"3f012d40", -- a1bc
		x"ffea4eba", -- a1c0
		x"ea22202e", -- a1c4
		x"ffea801f", -- a1c8
		x"67ca558f", -- a1cc
		x"2f2efffa", -- a1d0
		x"206effee", -- a1d4
		x"70001028", -- a1d8
		x"00023f00", -- a1dc
		x"4ebaea04", -- a1e0
		x"4a1f6700", -- a1e4
		x"01b01d7c", -- a1e8
		x"0001ffff", -- a1ec
		x"4a2e0008", -- a1f0
		x"67000032", -- a1f4
		x"206efff2", -- a1f8
		x"226effee", -- a1fc
		x"70001029", -- a200
		x"00023200", -- a204
		x"e841e349", -- a208
		x"0240000f", -- a20c
		x"45e802fc", -- a210
		x"24321000", -- a214
		x"e1aa701f", -- a218
		x"e0aa4a82", -- a21c
		x"67000006", -- a220
		x"422effff", -- a224
		x"4a2effff", -- a228
		x"6700016a", -- a22c
		x"206efff2", -- a230
		x"08280003", -- a234
		x"005c56c0", -- a238
		x"44004a00", -- a23c
		x"6600010c", -- a240
		x"2d6efff6", -- a244
		x"ffea2f2d", -- a248
		x"fff62f0e", -- a24c
		x"487a00ea", -- a250
		x"2b4ffff6", -- a254
		x"42a80092", -- a258
		x"42a80096", -- a25c
		x"08e80003", -- a260
		x"005c226e", -- a264
		x"fffa237c", -- a268
		x"00001388", -- a26c
		x"0004226e", -- a270
		x"ffee7000", -- a274
		x"10290002", -- a278
		x"2f002f3c", -- a27c
		x"000000ff", -- a280
		x"4ebaf26a", -- a284
		x"206effee", -- a288
		x"70001028", -- a28c
		x"00022f00", -- a290
		x"2f3c0000", -- a294
		x"00ff7000", -- a298
		x"10280001", -- a29c
		x"2f004eba", -- a2a0
		x"f3de206e", -- a2a4
		x"fff2226e", -- a2a8
		x"ffea7000", -- a2ac
		x"10290008", -- a2b0
		x"3200e841", -- a2b4
		x"e3490240", -- a2b8
		x"000f45e8", -- a2bc
		x"00927401", -- a2c0
		x"4400d03c", -- a2c4
		x"001fe1aa", -- a2c8
		x"4682c5b2", -- a2cc
		x"10007401", -- a2d0
		x"76001602", -- a2d4
		x"e1ab87b2", -- a2d8
		x"1000206e", -- a2dc
		x"ffee7000", -- a2e0
		x"10280002", -- a2e4
		x"2f002f3c", -- a2e8
		x"00000016", -- a2ec
		x"4ebaeb6e", -- a2f0
		x"206efff2", -- a2f4
		x"226effea", -- a2f8
		x"70001029", -- a2fc
		x"00083200", -- a300
		x"e841e349", -- a304
		x"0240000f", -- a308
		x"45e80092", -- a30c
		x"74014400", -- a310
		x"d03c001f", -- a314
		x"e1aa4682", -- a318
		x"c5b21000", -- a31c
		x"74017600", -- a320
		x"1602e1ab", -- a324
		x"87b21000", -- a328
		x"60b02b6f", -- a32c
		x"0008fff6", -- a330
		x"defc000c", -- a334
		x"4efa0014", -- a338
		x"2c5f2b5f", -- a33c
		x"fff67001", -- a340
		x"b06dfffe", -- a344
		x"67000004", -- a348
		x"4e4a206e", -- a34c
		x"fff22028", -- a350
		x"005eb0ba", -- a354
		x"e85e56c0", -- a358
		x"226effee", -- a35c
		x"72001229", -- a360
		x"00033401", -- a364
		x"e842e34a", -- a368
		x"0241000f", -- a36c
		x"45e80092", -- a370
		x"26322000", -- a374
		x"e3ab721f", -- a378
		x"e2abc003", -- a37c
		x"67000016", -- a380
		x"246e000e", -- a384
		x"24a8005e", -- a388
		x"558f4eba", -- a38c
		x"f35c206e", -- a390
		x"000a109f", -- a394
		x"6000fc60", -- a398
		x"206e000a", -- a39c
		x"1d500016", -- a3a0
		x"2b6f0008", -- a3a4
		x"fff6defc", -- a3a8
		x"000c4efa", -- a3ac
		x"00262c5f", -- a3b0
		x"2b5ffff6", -- a3b4
		x"422e0016", -- a3b8
		x"302dfffe", -- a3bc
		x"48c02f00", -- a3c0
		x"487a001a", -- a3c4
		x"4ebaddea", -- a3c8
		x"4a1f6600", -- a3cc
		x"00064eba", -- a3d0
		x"be744e5e", -- a3d4
		x"205fdefc", -- a3d8
		x"000e4ed0", -- a3dc
		x"00026000", -- a3e0
		x"00004e56", -- a3e4
		x"fff62f2d", -- a3e8
		x"fff62f0e", -- a3ec
		x"487a0038", -- a3f0
		x"2b4ffff6", -- a3f4
		x"3d7ce942", -- a3f8
		x"fff6558f", -- a3fc
		x"2f2e0008", -- a400
		x"486efff8", -- a404
		x"486efffc", -- a408
		x"486efff6", -- a40c
		x"4ebaf4a6", -- a410
		x"1d5f000c", -- a414
		x"4ebaf956", -- a418
		x"2b6f0008", -- a41c
		x"fff6defc", -- a420
		x"000c4efa", -- a424
		x"00102c5f", -- a428
		x"2b5ffff6", -- a42c
		x"422e000c", -- a430
		x"4ebabe12", -- a434
		x"4e5e2e9f", -- a438
		x"4e754e75", -- a43c
		x"241f40e7", -- a440
		x"2f02342f", -- a444
		x"0004c47c", -- a448
		x"f8ff847c", -- a44c
		x"060046c2", -- a450
		x"08380001", -- a454
		x"feda6622", -- a458
		x"2f3c000f", -- a45c
		x"42404857", -- a460
		x"4eb8521e", -- a464
		x"241f4a2b", -- a468
		x"00046a3a", -- a46c
		x"2f024857", -- a470
		x"4eb8523e", -- a474
		x"6aee588f", -- a478
		x"6010243c", -- a47c
		x"0002673c", -- a480
		x"4a2b0004", -- a484
		x"6a205382", -- a488
		x"66f646ef", -- a48c
		x"00046000", -- a490
		x"008c1740", -- a494
		x"000446ef", -- a498
		x"00043f6f", -- a49c
		x"00020004", -- a4a0
		x"3f570002", -- a4a4
		x"548f4e75", -- a4a8
		x"205f265f", -- a4ac
		x"524b2f08", -- a4b0
		x"422b400c", -- a4b4
		x"177c0080", -- a4b8
		x"00006180", -- a4bc
		x"61d451ef", -- a4c0
		x"00044a2b", -- a4c4
		x"400c6604", -- a4c8
		x"50ef0004", -- a4cc
		x"4e757a04", -- a4d0
		x"60027a24", -- a4d4
		x"45f80006", -- a4d8
		x"4284090b", -- a4dc
		x"4008ee5c", -- a4e0
		x"d88b2244", -- a4e4
		x"4284d3ca", -- a4e8
		x"09090000", -- a4ec
		x"ee5cd88b", -- a4f0
		x"d8852444", -- a4f4
		x"4e7543f8", -- a4f8
		x"00106004", -- a4fc
		x"43f80000", -- a500
		x"d3ca4285", -- a504
		x"0b090004", -- a508
		x"e05d4284", -- a50c
		x"09090000", -- a510
		x"ee5cd88b", -- a514
		x"2244d885", -- a518
		x"d8854e75", -- a51c
		x"70056002", -- a520
		x"70013b40", -- a524
		x"fffe4e4a", -- a528
		x"61cc4280", -- a52c
		x"4281030a", -- a530
		x"000c6100", -- a534
		x"ff08010a", -- a538
		x"0018050a", -- a53c
		x"00086100", -- a540
		x"ff52b242", -- a544
		x"670aee59", -- a548
		x"d28b2041", -- a54c
		x"01080000", -- a550
		x"e058030a", -- a554
		x"001ce059", -- a558
		x"90416c02", -- a55c
		x"d0454e75", -- a560
		x"619a4280", -- a564
		x"010a000c", -- a568
		x"ee58d08b", -- a56c
		x"2040d07c", -- a570
		x"0008b840", -- a574
		x"66023009", -- a578
		x"08800000", -- a57c
		x"ef586100", -- a580
		x"febc018a", -- a584
		x"000c6100", -- a588
		x"ff0a4e75", -- a58c
		x"619a2600", -- a590
		x"48e70020", -- a594
		x"4280010a", -- a598
		x"001cee58", -- a59c
		x"d08b2440", -- a5a0
		x"90844480", -- a5a4
		x"c0bc0000", -- a5a8
		x"fffee258", -- a5ac
		x"b6806e02", -- a5b0
		x"2003242c", -- a5b4
		x"000eb480", -- a5b8
		x"6e022002", -- a5bc
		x"26006738", -- a5c0
		x"5340206c", -- a5c4
		x"000a10d2", -- a5c8
		x"544a51c8", -- a5cc
		x"fffa9483", -- a5d0
		x"2942000e", -- a5d4
		x"2948000a", -- a5d8
		x"220ab88a", -- a5dc
		x"66022209", -- a5e0
		x"08810000", -- a5e4
		x"ef594cdf", -- a5e8
		x"04006100", -- a5ec
		x"fe50038a", -- a5f0
		x"001c6100", -- a5f4
		x"fe9e4e75", -- a5f8
		x"4cdf0400", -- a5fc
		x"4e756100", -- a600
		x"fef66100", -- a604
		x"fe38070a", -- a608
		x"0018030a", -- a60c
		x"00086100", -- a610
		x"fe824282", -- a614
		x"4280050a", -- a618
		x"000cb441", -- a61c
		x"660c050a", -- a620
		x"001cb443", -- a624
		x"67025200", -- a628
		x"4e755400", -- a62c
		x"60f06100", -- a630
		x"fe0c050a", -- a634
		x"00086100", -- a638
		x"fe5a4280", -- a63c
		x"010a000c", -- a640
		x"b4406716", -- a644
		x"ee58d08b", -- a648
		x"20400108", -- a64c
		x"00004285", -- a650
		x"050a001c", -- a654
		x"b44057c0", -- a658
		x"4e754280", -- a65c
		x"4e75205f", -- a660
		x"221f225f", -- a664
		x"285f4850", -- a668
		x"266c0000", -- a66c
		x"528b2949", -- a670
		x"000a2941", -- a674
		x"000e296c", -- a678
		x"00040016", -- a67c
		x"08380001", -- a680
		x"feda6612", -- a684
		x"486c0016", -- a688
		x"4eb851f4", -- a68c
		x"486c0016", -- a690
		x"4eb8521e", -- a694
		x"6008297c", -- a698
		x"00000007", -- a69c
		x"001a6100", -- a6a0
		x"fe2e6746", -- a6a4
		x"4aac000e", -- a6a8
		x"67406100", -- a6ac
		x"01b04a2b", -- a6b0
		x"400c6600", -- a6b4
		x"fe6c0838", -- a6b8
		x"0001feda", -- a6bc
		x"660e486c", -- a6c0
		x"00164eb8", -- a6c4
		x"523e6adc", -- a6c8
		x"6000fe56", -- a6cc
		x"53ac001a", -- a6d0
		x"66d2297c", -- a6d4
		x"00000007", -- a6d8
		x"001a4aac", -- a6dc
		x"001667c4", -- a6e0
		x"53ac0016", -- a6e4
		x"6700fe3a", -- a6e8
		x"60ba4e75", -- a6ec
		x"205f245f", -- a6f0
		x"225f285f", -- a6f4
		x"4850266c", -- a6f8
		x"0000528b", -- a6fc
		x"2949000a", -- a700
		x"296c0004", -- a704
		x"00160838", -- a708
		x"0001feda", -- a70c
		x"6612486c", -- a710
		x"00164eb8", -- a714
		x"51f4486c", -- a718
		x"00164eb8", -- a71c
		x"521e6008", -- a720
		x"297c0000", -- a724
		x"0006001a", -- a728
		x"2952000e", -- a72c
		x"2f0a6006", -- a730
		x"4aac000e", -- a734
		x"675c6100", -- a738
		x"fd9a4a2b", -- a73c
		x"400c6600", -- a740
		x"fde00838", -- a744
		x"0001feda", -- a748
		x"660c486c", -- a74c
		x"00164eb8", -- a750
		x"523e6a2a", -- a754
		x"601a53ac", -- a758
		x"001a6622", -- a75c
		x"297c0000", -- a760
		x"0006001a", -- a764
		x"4aac0016", -- a768
		x"671453ac", -- a76c
		x"0016660e", -- a770
		x"205f2010", -- a774
		x"90ac000e", -- a778
		x"20806000", -- a77c
		x"fda46100", -- a780
		x"fe7e4a00", -- a784
		x"67aa6100", -- a788
		x"fea64a00", -- a78c
		x"67106100", -- a790
		x"fdd0205f", -- a794
		x"201090ac", -- a798
		x"000e2080", -- a79c
		x"4e754aac", -- a7a0
		x"000e67ee", -- a7a4
		x"6100fde6", -- a7a8
		x"6086205f", -- a7ac
		x"285f4850", -- a7b0
		x"266c0000", -- a7b4
		x"528b6100", -- a7b8
		x"fd16296c", -- a7bc
		x"00040012", -- a7c0
		x"08380001", -- a7c4
		x"feda6612", -- a7c8
		x"486c0012", -- a7cc
		x"4eb851f4", -- a7d0
		x"486c0012", -- a7d4
		x"4eb8521e", -- a7d8
		x"6008297c", -- a7dc
		x"0000000b", -- a7e0
		x"001e6100", -- a7e4
		x"01864a00", -- a7e8
		x"663c4a2b", -- a7ec
		x"400c6600", -- a7f0
		x"fd300838", -- a7f4
		x"0001feda", -- a7f8
		x"660e486c", -- a7fc
		x"00124eb8", -- a800
		x"523e6ade", -- a804
		x"6000fd1a", -- a808
		x"53ac001e", -- a80c
		x"66d4297c", -- a810
		x"0000000b", -- a814
		x"001e4aac", -- a818
		x"001267c6", -- a81c
		x"53ac0012", -- a820
		x"66c06000", -- a824
		x"fcfc4e75", -- a828
		x"42804283", -- a82c
		x"010a0008", -- a830
		x"6100fc0a", -- a834
		x"070a000c", -- a838
		x"60104280", -- a83c
		x"4283010a", -- a840
		x"00186100", -- a844
		x"fbf8070a", -- a848
		x"001c6100", -- a84c
		x"fc46e058", -- a850
		x"e05b9640", -- a854
		x"53436c02", -- a858
		x"d6454e75", -- a85c
		x"6100fc98", -- a860
		x"61d82200", -- a864
		x"20040280", -- a868
		x"0000fffe", -- a86c
		x"e2809081", -- a870
		x"b6806e02", -- a874
		x"2003242c", -- a878
		x"000eb480", -- a87c
		x"6e022002", -- a880
		x"26006740", -- a884
		x"5340206c", -- a888
		x"000ae349", -- a88c
		x"d28b48e7", -- a890
		x"00402241", -- a894
		x"12985449", -- a898
		x"51c8fffa", -- a89c
		x"94832942", -- a8a0
		x"000e2948", -- a8a4
		x"000a2209", -- a8a8
		x"4cdf0200", -- a8ac
		x"b8816602", -- a8b0
		x"22090881", -- a8b4
		x"0000ef59", -- a8b8
		x"6100fb82", -- a8bc
		x"038a0018", -- a8c0
		x"6100fbd0", -- a8c4
		x"4e756100", -- a8c8
		x"fc066100", -- a8cc
		x"fc30296c", -- a8d0
		x"00040012", -- a8d4
		x"08380001", -- a8d8
		x"feda6612", -- a8dc
		x"486c0012", -- a8e0
		x"4eb851f4", -- a8e4
		x"486c0012", -- a8e8
		x"4eb8521e", -- a8ec
		x"6008297c", -- a8f0
		x"0000000b", -- a8f4
		x"001e6100", -- a8f8
		x"ff300c83", -- a8fc
		x"00000004", -- a900
		x"6c340838", -- a904
		x"0001feda", -- a908
		x"660e486c", -- a90c
		x"00124eb8", -- a910
		x"523e6ae2", -- a914
		x"6000fc0a", -- a918
		x"53ac001e", -- a91c
		x"66d8297c", -- a920
		x"0000000b", -- a924
		x"001e4aac", -- a928
		x"001267ca", -- a92c
		x"53ac0012", -- a930
		x"66c46000", -- a934
		x"fbece348", -- a938
		x"d08b2040", -- a93c
		x"010a0018", -- a940
		x"01880000", -- a944
		x"302c0008", -- a948
		x"01880004", -- a94c
		x"50882208", -- a950
		x"b8816602", -- a954
		x"22090881", -- a958
		x"0000ef59", -- a95c
		x"6100fade", -- a960
		x"038a0008", -- a964
		x"6100fb2c", -- a968
		x"4e757204", -- a96c
		x"4280102a", -- a970
		x"fffc6714", -- a974
		x"22006100", -- a978
		x"fb7e6100", -- a97c
		x"febeb681", -- a980
		x"6c044280", -- a984
		x"4e757208", -- a988
		x"6100fb72", -- a98c
		x"6100fe9a", -- a990
		x"b6816dee", -- a994
		x"397c0500", -- a998
		x"00086100", -- a99c
		x"ff2a7001", -- a9a0
		x"4e75ffff", -- a9a4
		x"5d06ee1b", -- a9a8
		x"ffff4e75", -- a9ac
		x"611601d0", -- a9b0
		x"4ed16110", -- a9b4
		x"01904ed1", -- a9b8
		x"610a0110", -- a9bc
		x"56c04400", -- a9c0
		x"1e804ed1", -- a9c4
		x"245f225f", -- a9c8
		x"301f305f", -- a9cc
		x"d1df4ed2", -- a9d0
		x"205f201f", -- a9d4
		x"c09f2e80", -- a9d8
		x"4ed0205f", -- a9dc
		x"201f4680", -- a9e0
		x"2e804ed0", -- a9e4
		x"2078fed4", -- a9e8
		x"10280060", -- a9ec
		x"488048c0", -- a9f0
		x"6b1cb03c", -- a9f4
		x"00076610", -- a9f8
		x"08380005", -- a9fc
		x"fed26608", -- aa00
		x"203c0047", -- aa04
		x"80006006", -- aa08
		x"807c0060", -- aa0c
		x"4840205f", -- aa10
		x"2e804ed0", -- aa14
		x"598f61cc", -- aa18
		x"225f6b20", -- aa1c
		x"7020b3fc", -- aa20
		x"00478000", -- aa24
		x"67167000", -- aa28
		x"2478fed4", -- aa2c
		x"122a0060", -- aa30
		x"6100d5c4", -- aa34
		x"6706707f", -- aa38
		x"c0290001", -- aa3c
		x"205f3e80", -- aa40
		x"4ed0205f", -- aa44
		x"225f245f", -- aa48
		x"72097020", -- aa4c
		x"b0311000", -- aa50
		x"56c9fffa", -- aa54
		x"52412649", -- aa58
		x"1601284a", -- aa5c
		x"181c5304", -- aa60
		x"650e101c", -- aa64
		x"670e5303", -- aa68
		x"651cb01b", -- aa6c
		x"661860ee", -- aa70
		x"53036412", -- aa74
		x"14c15301", -- aa78
		x"650614d9", -- aa7c
		x"51c9fffc", -- aa80
		x"1ebc0001", -- aa84
		x"4ed051d7", -- aa88
		x"4ed00838", -- aa8c
		x"0001feda", -- aa90
		x"6700a7d8", -- aa94
		x"2f2f0004", -- aa98
		x"2f6f0004", -- aa9c
		x"00082f40", -- aaa0
		x"0004201f", -- aaa4
		x"51c8fffe", -- aaa8
		x"42405380", -- aaac
		x"64f6201f", -- aab0
		x"4e75e200", -- aab4
		x"0000e200", -- aab8
		x"15000000", -- aabc
		x"4e56fff4", -- aac0
		x"2d7c0000", -- aac4
		x"03e8fffc", -- aac8
		x"2d6e0008", -- aacc
		x"fff8206e", -- aad0
		x"fff82d68", -- aad4
		x"0002fff4", -- aad8
		x"206efff4", -- aadc
		x"226e000c", -- aae0
		x"32a84000", -- aae4
		x"53aefffc", -- aae8
		x"4aaefffc", -- aaec
		x"5fc00828", -- aaf0
		x"00020003", -- aaf4
		x"56c14401", -- aaf8
		x"800167dc", -- aafc
		x"08280002", -- ab00
		x"000356c0", -- ab04
		x"44004a00", -- ab08
		x"66000018", -- ab0c
		x"226efff8", -- ab10
		x"32bc0002", -- ab14
		x"117c0001", -- ab18
		x"00013b7c", -- ab1c
		x"0005fffe", -- ab20
		x"4e4a4e5e", -- ab24
		x"205f504f", -- ab28
		x"4ed00000", -- ab2c
		x"4e56fff4", -- ab30
		x"2d7c0000", -- ab34
		x"03e8fffc", -- ab38
		x"2d6e000c", -- ab3c
		x"fff8206e", -- ab40
		x"fff82d68", -- ab44
		x"0002fff4", -- ab48
		x"206efff4", -- ab4c
		x"316e000a", -- ab50
		x"400053ae", -- ab54
		x"fffc4aae", -- ab58
		x"fffc5fc0", -- ab5c
		x"08280002", -- ab60
		x"000356c1", -- ab64
		x"44018001", -- ab68
		x"67de0828", -- ab6c
		x"00020003", -- ab70
		x"56c04400", -- ab74
		x"4a006600", -- ab78
		x"0018226e", -- ab7c
		x"fff832bc", -- ab80
		x"0002117c", -- ab84
		x"00010001", -- ab88
		x"3b7c0005", -- ab8c
		x"fffe4e4a", -- ab90
		x"4e5e205f", -- ab94
		x"504f4ed0", -- ab98
		x"00004e56", -- ab9c
		x"ffde2d6e", -- aba0
		x"0008ffee", -- aba4
		x"206effee", -- aba8
		x"2d680002", -- abac
		x"ffea226e", -- abb0
		x"ffea137c", -- abb4
		x"ff010001", -- abb8
		x"d3fc0000", -- abbc
		x"800043d1", -- abc0
		x"2d49fffc", -- abc4
		x"226effea", -- abc8
		x"337c0001", -- abcc
		x"4002302e", -- abd0
		x"fffe3340", -- abd4
		x"4000337c", -- abd8
		x"00024002", -- abdc
		x"102efffd", -- abe0
		x"024000ff", -- abe4
		x"33404000", -- abe8
		x"337c0003", -- abec
		x"4002337c", -- abf0
		x"00044000", -- abf4
		x"d3fc0000", -- abf8
		x"800043d1", -- abfc
		x"2d49ffe6", -- ac00
		x"226effe6", -- ac04
		x"2d49ffe2", -- ac08
		x"246effe2", -- ac0c
		x"34bc0000", -- ac10
		x"08920007", -- ac14
		x"15680009", -- ac18
		x"00021568", -- ac1c
		x"00080003", -- ac20
		x"1568000b", -- ac24
		x"00041568", -- ac28
		x"000a0005", -- ac2c
		x"1568000d", -- ac30
		x"00061568", -- ac34
		x"000c0007", -- ac38
		x"4cb91b00", -- ac3c
		x"0000dcee", -- ac40
		x"48aa1b00", -- ac44
		x"0008206e", -- ac48
		x"ffe643e8", -- ac4c
		x"00182d49", -- ac50
		x"fffc302e", -- ac54
		x"fffe3540", -- ac58
		x"0010156e", -- ac5c
		x"fffd0013", -- ac60
		x"022aff1f", -- ac64
		x"00127004", -- ac68
		x"eb88812a", -- ac6c
		x"0012022a", -- ac70
		x"00e00012", -- ac74
		x"7000812a", -- ac78
		x"001243e8", -- ac7c
		x"00982d49", -- ac80
		x"fffc302e", -- ac84
		x"fffe3540", -- ac88
		x"0014156e", -- ac8c
		x"fffd0017", -- ac90
		x"022aff1f", -- ac94
		x"00167000", -- ac98
		x"eb88812a", -- ac9c
		x"0016022a", -- aca0
		x"00e00016", -- aca4
		x"7000812a", -- aca8
		x"0016426e", -- acac
		x"fff6526e", -- acb0
		x"fff6206e", -- acb4
		x"ffe6302e", -- acb8
		x"fff648c0", -- acbc
		x"e78043f0", -- acc0
		x"08102d49", -- acc4
		x"ffde302e", -- acc8
		x"fff6c1fc", -- accc
		x"03c443e8", -- acd0
		x"fcdc43f1", -- acd4
		x"08002d49", -- acd8
		x"fffc226e", -- acdc
		x"ffde302e", -- ace0
		x"fffe3280", -- ace4
		x"136efffd", -- ace8
		x"0003137c", -- acec
		x"ff800002", -- acf0
		x"337cfc3c", -- acf4
		x"00044269", -- acf8
		x"00060c6e", -- acfc
		x"0010fff6", -- ad00
		x"6dac206e", -- ad04
		x"ffee317c", -- ad08
		x"00010006", -- ad0c
		x"226effe6", -- ad10
		x"137cff00", -- ad14
		x"009a246e", -- ad18
		x"ffea357c", -- ad1c
		x"00004002", -- ad20
		x"35790000", -- ad24
		x"dcec4000", -- ad28
		x"2d7c0000", -- ad2c
		x"7530fff8", -- ad30
		x"486efff8", -- ad34
		x"4ebaa4e4", -- ad38
		x"422efff5", -- ad3c
		x"2f2dfff6", -- ad40
		x"2f0e487a", -- ad44
		x"00c82b4f", -- ad48
		x"fff6206e", -- ad4c
		x"ffea0828", -- ad50
		x"00060003", -- ad54
		x"56c04400", -- ad58
		x"4a006700", -- ad5c
		x"007e486e", -- ad60
		x"ffe02f2e", -- ad64
		x"00084eba", -- ad68
		x"fd543d6e", -- ad6c
		x"ffe0fff2", -- ad70
		x"082e0000", -- ad74
		x"fff256c0", -- ad78
		x"44004a00", -- ad7c
		x"6700005c", -- ad80
		x"082e0000", -- ad84
		x"fff356c0", -- ad88
		x"4400082e", -- ad8c
		x"0001fff3", -- ad90
		x"56c14401", -- ad94
		x"c200082e", -- ad98
		x"0004fff3", -- ad9c
		x"56c04400", -- ada0
		x"c001082e", -- ada4
		x"0006fff3", -- ada8
		x"56c14401", -- adac
		x"c2006600", -- adb0
		x"000a3b7c", -- adb4
		x"0005fffe", -- adb8
		x"4e4a2f2e", -- adbc
		x"00087000", -- adc0
		x"30390000", -- adc4
		x"dcea2f00", -- adc8
		x"4ebafd62", -- adcc
		x"1d7cfd01", -- add0
		x"fff5206e", -- add4
		x"ffee30bc", -- add8
		x"0005558f", -- addc
		x"486efff8", -- ade0
		x"4ebaa472", -- ade4
		x"101f802e", -- ade8
		x"fff56700", -- adec
		x"ff5e4a2e", -- adf0
		x"fff56600", -- adf4
		x"000a3b7c", -- adf8
		x"0005fffe", -- adfc
		x"4e4a2b6f", -- ae00
		x"0008fff6", -- ae04
		x"defc000c", -- ae08
		x"4efa003a", -- ae0c
		x"2c5f2b5f", -- ae10
		x"fff67005", -- ae14
		x"b06dfffe", -- ae18
		x"66000028", -- ae1c
		x"206effee", -- ae20
		x"7002b050", -- ae24
		x"67000006", -- ae28
		x"30bc0001", -- ae2c
		x"206effea", -- ae30
		x"117cff01", -- ae34
		x"00013b7c", -- ae38
		x"0005fffe", -- ae3c
		x"4e4a6000", -- ae40
		x"00044e4a", -- ae44
		x"4e5e2e9f", -- ae48
		x"4e750000", -- ae4c
		x"4e56fff8", -- ae50
		x"2079ffff", -- ae54
		x"fed4302e", -- ae58
		x"00083200", -- ae5c
		x"e841e349", -- ae60
		x"0240000f", -- ae64
		x"41e800dc", -- ae68
		x"24301000", -- ae6c
		x"e1aa701f", -- ae70
		x"e0aa4a82", -- ae74
		x"6700006a", -- ae78
		x"2d6e000a", -- ae7c
		x"fffc2f3c", -- ae80
		x"00010000", -- ae84
		x"7060d06e", -- ae88
		x"000848c0", -- ae8c
		x"2f004eba", -- ae90
		x"d31c206e", -- ae94
		x"fffc215f", -- ae98
		x"00022d68", -- ae9c
		x"0002fff8", -- aea0
		x"226efff8", -- aea4
		x"10290001", -- aea8
		x"02800000", -- aeac
		x"007f7215", -- aeb0
		x"b2806600", -- aeb4
		x"00084250", -- aeb8
		x"6000000a", -- aebc
		x"3b7c0001", -- aec0
		x"fffe4e4a", -- aec4
		x"206efff8", -- aec8
		x"117cff01", -- aecc
		x"0001117c", -- aed0
		x"ff000003", -- aed4
		x"226efffc", -- aed8
		x"32bc0004", -- aedc
		x"6000000a", -- aee0
		x"3b7c0001", -- aee4
		x"fffe4e4a", -- aee8
		x"4e5e205f", -- aeec
		x"5c4f4ed0", -- aef0
		x"00004e56", -- aef4
		x"fff82f2d", -- aef8
		x"fff62f0e", -- aefc
		x"487a006c", -- af00
		x"2b4ffff6", -- af04
		x"2d6e000a", -- af08
		x"fffc2d79", -- af0c
		x"fffffed4", -- af10
		x"fff82f2e", -- af14
		x"000a206e", -- af18
		x"fff87000", -- af1c
		x"10280060", -- af20
		x"3f004eba", -- af24
		x"ff28558f", -- af28
		x"206efffc", -- af2c
		x"2f280002", -- af30
		x"48680008", -- af34
		x"4eba2850", -- af38
		x"4a1f6600", -- af3c
		x"000a3b7c", -- af40
		x"0005fffe", -- af44
		x"4e4a2f2e", -- af48
		x"000a4eba", -- af4c
		x"fc4e206e", -- af50
		x"fffc4268", -- af54
		x"00141d7c", -- af58
		x"0001000e", -- af5c
		x"2b6f0008", -- af60
		x"fff6defc", -- af64
		x"000c4efa", -- af68
		x"00242c5f", -- af6c
		x"2b5ffff6", -- af70
		x"422e000e", -- af74
		x"302dfffe", -- af78
		x"48c02f00", -- af7c
		x"487a0016", -- af80
		x"4ebad22e", -- af84
		x"4a1f6600", -- af88
		x"00044e4a", -- af8c
		x"4e5e205f", -- af90
		x"5c4f4ed0", -- af94
		x"00024400", -- af98
		x"00004e56", -- af9c
		x"fff4206e", -- afa0
		x"000a2068", -- afa4
		x"0002d1fc", -- afa8
		x"00008000", -- afac
		x"41d02d48", -- afb0
		x"fff80c6e", -- afb4
		x"03200008", -- afb8
		x"6f00000a", -- afbc
		x"3b7c0006", -- afc0
		x"fffe4e4a", -- afc4
		x"206efff8", -- afc8
		x"43e83ce0", -- afcc
		x"2d49fffc", -- afd0
		x"43e80098", -- afd4
		x"2d49fff4", -- afd8
		x"302e0008", -- afdc
		x"4440226e", -- afe0
		x"fff43340", -- afe4
		x"0004337c", -- afe8
		x"00000006", -- afec
		x"302efffe", -- aff0
		x"3280136e", -- aff4
		x"fffd0003", -- aff8
		x"4e5e205f", -- affc
		x"5c4f4ed0", -- b000
		x"00004e56", -- b004
		x"0000558f", -- b008
		x"2f2e0008", -- b00c
		x"2079ffff", -- b010
		x"fed47000", -- b014
		x"10280060", -- b018
		x"3f004eba", -- b01c
		x"fed64a1f", -- b020
		x"6600000a", -- b024
		x"3b7c0005", -- b028
		x"fffe4e4a", -- b02c
		x"4e5e2e9f", -- b030
		x"4e750000", -- b034
		x"4e56fff2", -- b038
		x"2d6e0008", -- b03c
		x"fff8206e", -- b040
		x"fff82d68", -- b044
		x"0002fff4", -- b048
		x"226efff4", -- b04c
		x"08290001", -- b050
		x"000356c0", -- b054
		x"44004a00", -- b058
		x"67000012", -- b05c
		x"2f2e0008", -- b060
		x"4ebaffa0", -- b064
		x"3b7cffff", -- b068
		x"fffe4e4a", -- b06c
		x"486efff2", -- b070
		x"2f2e0008", -- b074
		x"4ebafa46", -- b078
		x"3d6efff2", -- b07c
		x"fffe206e", -- b080
		x"000c30ae", -- b084
		x"fffe2f2e", -- b088
		x"0008558f", -- b08c
		x"3f2efffe", -- b090
		x"3f390000", -- b094
		x"dce64eba", -- b098
		x"26b6301f", -- b09c
		x"48c02f00", -- b0a0
		x"4ebafa8a", -- b0a4
		x"082e0003", -- b0a8
		x"fffe56c0", -- b0ac
		x"4400082e", -- b0b0
		x"0006fffe", -- b0b4
		x"56c14401", -- b0b8
		x"8200082e", -- b0bc
		x"0007fffe", -- b0c0
		x"56c04400", -- b0c4
		x"c2006700", -- b0c8
		x"0014206e", -- b0cc
		x"fff4117c", -- b0d0
		x"ff010001", -- b0d4
		x"3b7c0005", -- b0d8
		x"fffe4e4a", -- b0dc
		x"4e5e205f", -- b0e0
		x"504f4ed0", -- b0e4
		x"00004e56", -- b0e8
		x"fff8422e", -- b0ec
		x"000c2d6e", -- b0f0
		x"0008fffc", -- b0f4
		x"206efffc", -- b0f8
		x"22680002", -- b0fc
		x"d3fc0000", -- b100
		x"809843d1", -- b104
		x"2d49fff8", -- b108
		x"226efff8", -- b10c
		x"08290007", -- b110
		x"000256c0", -- b114
		x"44004a00", -- b118
		x"6600005c", -- b11c
		x"08290006", -- b120
		x"000656c0", -- b124
		x"44000829", -- b128
		x"00070006", -- b12c
		x"56c14401", -- b130
		x"82006700", -- b134
		x"00202468", -- b138
		x"0002157c", -- b13c
		x"00010001", -- b140
		x"2f2e0008", -- b144
		x"4ebafebc", -- b148
		x"3b7cffff", -- b14c
		x"fffe4e4a", -- b150
		x"60000024", -- b154
		x"1d7c0001", -- b158
		x"000c206e", -- b15c
		x"fff80828", -- b160
		x"00060002", -- b164
		x"56c04400", -- b168
		x"4a006700", -- b16c
		x"000a3b7c", -- b170
		x"fffefffe", -- b174
		x"4e4a4e5e", -- b178
		x"2e9f4e75", -- b17c
		x"00004e56", -- b180
		x"ffea426e", -- b184
		x"fffe2d6e", -- b188
		x"0010fff6", -- b18c
		x"206efff6", -- b190
		x"22680002", -- b194
		x"d3fc0000", -- b198
		x"800043d1", -- b19c
		x"2d49fff2", -- b1a0
		x"226efff2", -- b1a4
		x"30280006", -- b1a8
		x"48c0e780", -- b1ac
		x"45f10810", -- b1b0
		x"2d4affee", -- b1b4
		x"246effee", -- b1b8
		x"082a0007", -- b1bc
		x"000256c0", -- b1c0
		x"44004a00", -- b1c4
		x"6700000c", -- b1c8
		x"3d7c0001", -- b1cc
		x"00146000", -- b1d0
		x"00f2206e", -- b1d4
		x"ffee0828", -- b1d8
		x"00010002", -- b1dc
		x"56c04400", -- b1e0
		x"4a006600", -- b1e4
		x"000c3d7c", -- b1e8
		x"00020014", -- b1ec
		x"600000d4", -- b1f0
		x"206efff6", -- b1f4
		x"3d680006", -- b1f8
		x"fffa3d7c", -- b1fc
		x"0003fffc", -- b200
		x"206efff2", -- b204
		x"302efffa", -- b208
		x"48c0e780", -- b20c
		x"43f00810", -- b210
		x"2d49ffea", -- b214
		x"226effea", -- b218
		x"08290007", -- b21c
		x"000256c0", -- b220
		x"44004a00", -- b224
		x"6700000c", -- b228
		x"3d7c0001", -- b22c
		x"fffc6000", -- b230
		x"0082558f", -- b234
		x"3f2efffe", -- b238
		x"206effea", -- b23c
		x"70001028", -- b240
		x"00023f00", -- b244
		x"4eba2512", -- b248
		x"3d5ffffe", -- b24c
		x"206effea", -- b250
		x"08280006", -- b254
		x"000256c0", -- b258
		x"44004a00", -- b25c
		x"6700000c", -- b260
		x"3d7c0002", -- b264
		x"fffc6000", -- b268
		x"004a206e", -- b26c
		x"ffea0828", -- b270
		x"00000002", -- b274
		x"56c04400", -- b278
		x"4a006700", -- b27c
		x"0012226e", -- b280
		x"000832a8", -- b284
		x"0006426e", -- b288
		x"fffc6000", -- b28c
		x"0026302e", -- b290
		x"fffa0240", -- b294
		x"000f5240", -- b298
		x"3d40fffa", -- b29c
		x"206efff6", -- b2a0
		x"302efffa", -- b2a4
		x"b0680006", -- b2a8
		x"66000008", -- b2ac
		x"3d7c0002", -- b2b0
		x"fffc7003", -- b2b4
		x"b06efffc", -- b2b8
		x"6700ff46", -- b2bc
		x"3d6efffc", -- b2c0
		x"0014206e", -- b2c4
		x"000c10ae", -- b2c8
		x"fffe4e5e", -- b2cc
		x"205fdefc", -- b2d0
		x"000c4ed0", -- b2d4
		x"00004e56", -- b2d8
		x"fff42d6e", -- b2dc
		x"0008fffc", -- b2e0
		x"206efffc", -- b2e4
		x"22680002", -- b2e8
		x"d3fc0000", -- b2ec
		x"800043d1", -- b2f0
		x"2d49fff8", -- b2f4
		x"206efff8", -- b2f8
		x"226efffc", -- b2fc
		x"30290006", -- b300
		x"48c0e780", -- b304
		x"45f00810", -- b308
		x"2d4afff4", -- b30c
		x"246efff4", -- b310
		x"426a0006", -- b314
		x"157c0080", -- b318
		x"00023029", -- b31c
		x"00060240", -- b320
		x"000f5240", -- b324
		x"33400006", -- b328
		x"30290006", -- b32c
		x"48c0e780", -- b330
		x"08300001", -- b334
		x"081256c0", -- b338
		x"44003229", -- b33c
		x"000648c1", -- b340
		x"e7810830", -- b344
		x"00071812", -- b348
		x"56c14401", -- b34c
		x"820067a4", -- b350
		x"4e5e2e9f", -- b354
		x"4e750000", -- b358
		x"4e56fff2", -- b35c
		x"2d6e0008", -- b360
		x"fffa206e", -- b364
		x"fffa2268", -- b368
		x"0002d3fc", -- b36c
		x"00008000", -- b370
		x"43d12d49", -- b374
		x"fff6206e", -- b378
		x"fff6226e", -- b37c
		x"fffa3029", -- b380
		x"000648c0", -- b384
		x"e78045f0", -- b388
		x"08102d4a", -- b38c
		x"fff2246e", -- b390
		x"fff2082a", -- b394
		x"00000002", -- b398
		x"56c04400", -- b39c
		x"082a0006", -- b3a0
		x"000256c1", -- b3a4
		x"44018200", -- b3a8
		x"02010001", -- b3ac
		x"1d41ffff", -- b3b0
		x"426a0006", -- b3b4
		x"157c0080", -- b3b8
		x"00023029", -- b3bc
		x"00060240", -- b3c0
		x"000f5240", -- b3c4
		x"33400006", -- b3c8
		x"4a2effff", -- b3cc
		x"67a84e5e", -- b3d0
		x"2e9f4e75", -- b3d4
		x"00004e56", -- b3d8
		x"ffe8422e", -- b3dc
		x"ffff422e", -- b3e0
		x"00102d6e", -- b3e4
		x"000cfff4", -- b3e8
		x"558f2f2e", -- b3ec
		x"000c486e", -- b3f0
		x"fffe486e", -- b3f4
		x"fffc4eba", -- b3f8
		x"fd863d5f", -- b3fc
		x"fffa302e", -- b400
		x"fffae340", -- b404
		x"323b0006", -- b408
		x"4efb1002", -- b40c
		x"0012014c", -- b410
		x"00062f2e", -- b414
		x"000c4eba", -- b418
		x"febe6000", -- b41c
		x"01420c6e", -- b420
		x"05eefffc", -- b424
		x"5ec07240", -- b428
		x"b26efffc", -- b42c
		x"5ec18200", -- b430
		x"6700000e", -- b434
		x"2f2e000c", -- b438
		x"4ebafe9c", -- b43c
		x"60000116", -- b440
		x"206efff4", -- b444
		x"22680002", -- b448
		x"d3fc0000", -- b44c
		x"800043d1", -- b450
		x"2d49fff0", -- b454
		x"226efff0", -- b458
		x"30280006", -- b45c
		x"48c0e780", -- b460
		x"45f10810", -- b464
		x"2d4affec", -- b468
		x"246e0008", -- b46c
		x"4292246e", -- b470
		x"ffec266e", -- b474
		x"00083012", -- b478
		x"37400002", -- b47c
		x"266e0008", -- b480
		x"176a0003", -- b484
		x"0001266e", -- b488
		x"00082d53", -- b48c
		x"ffe8266e", -- b490
		x"ffe80c6b", -- b494
		x"0640000c", -- b498
		x"54c01213", -- b49c
		x"c23c0601", -- b4a0
		x"80017203", -- b4a4
		x"b22b0010", -- b4a8
		x"56c18200", -- b4ac
		x"7000102b", -- b4b0
		x"000e0c40", -- b4b4
		x"00f856c0", -- b4b8
		x"80010c6b", -- b4bc
		x"06090014", -- b4c0
		x"56c18200", -- b4c4
		x"7000302b", -- b4c8
		x"000c740e", -- b4cc
		x"d0825880", -- b4d0
		x"342efffc", -- b4d4
		x"48c2b480", -- b4d8
		x"5dc08001", -- b4dc
		x"0200ff01", -- b4e0
		x"1d40fff9", -- b4e4
		x"4a2efff9", -- b4e8
		x"66000062", -- b4ec
		x"4cab1600", -- b4f0
		x"000648a8", -- b4f4
		x"1600000e", -- b4f8
		x"1d7c1601", -- b4fc
		x"00101d7c", -- b500
		x"1601ffff", -- b504
		x"226e0008", -- b508
		x"06910000", -- b50c
		x"00187000", -- b510
		x"302b000c", -- b514
		x"720ed081", -- b518
		x"72189081", -- b51c
		x"3140001e", -- b520
		x"7000302b", -- b524
		x"000c720e", -- b528
		x"d0813140", -- b52c
		x"00200c68", -- b530
		x"03c40020", -- b534
		x"6f000008", -- b538
		x"317c03c4", -- b53c
		x"0020206e", -- b540
		x"fff40468", -- b544
		x"00180020", -- b548
		x"6000000a", -- b54c
		x"2f2e000c", -- b550
		x"4ebafe06", -- b554
		x"60000008", -- b558
		x"1d7c0001", -- b55c
		x"ffff4a2e", -- b560
		x"ffff6700", -- b564
		x"fe844e5e", -- b568
		x"205f504f", -- b56c
		x"4ed00000", -- b570
		x"4e56ffee", -- b574
		x"206e0008", -- b578
		x"20680002", -- b57c
		x"d1fc0000", -- b580
		x"809a10bc", -- b584
		x"00832f2e", -- b588
		x"00087000", -- b58c
		x"30390000", -- b590
		x"dce42f00", -- b594
		x"4ebaf596", -- b598
		x"3d7c0003", -- b59c
		x"000c2d7c", -- b5a0
		x"003d0900", -- b5a4
		x"fffc486e", -- b5a8
		x"fffc4eba", -- b5ac
		x"9c6e2f2d", -- b5b0
		x"fff62f0e", -- b5b4
		x"487a00fc", -- b5b8
		x"2b4ffff6", -- b5bc
		x"2d6e0008", -- b5c0
		x"fff4206e", -- b5c4
		x"fff42d68", -- b5c8
		x"0002fff0", -- b5cc
		x"3d7c0001", -- b5d0
		x"fffa302e", -- b5d4
		x"fffa5340", -- b5d8
		x"e340323b", -- b5dc
		x"00064efb", -- b5e0
		x"10020006", -- b5e4
		x"00360058", -- b5e8
		x"206efff0", -- b5ec
		x"08280006", -- b5f0
		x"000356c0", -- b5f4
		x"44004a00", -- b5f8
		x"67000014", -- b5fc
		x"486effee", -- b600
		x"2f2e0008", -- b604
		x"4ebafa2e", -- b608
		x"3d6effee", -- b60c
		x"fff83d7c", -- b610
		x"0002fffa", -- b614
		x"60000086", -- b618
		x"558f2f2e", -- b61c
		x"00084eba", -- b620
		x"fac64a1f", -- b624
		x"6700000a", -- b628
		x"426efffa", -- b62c
		x"60000008", -- b630
		x"3d7c0003", -- b634
		x"fffa6000", -- b638
		x"0064206e", -- b63c
		x"fff00828", -- b640
		x"00060003", -- b644
		x"56c04400", -- b648
		x"4a006700", -- b64c
		x"002e486e", -- b650
		x"ffee2f2e", -- b654
		x"00084eba", -- b658
		x"f9dc3d6e", -- b65c
		x"ffeefff8", -- b660
		x"082e0001", -- b664
		x"fff856c0", -- b668
		x"44004a00", -- b66c
		x"67000008", -- b670
		x"3d7c0002", -- b674
		x"fffa6000", -- b678
		x"0024558f", -- b67c
		x"486efffc", -- b680
		x"4eba9bd2", -- b684
		x"4a1f6700", -- b688
		x"0014206e", -- b68c
		x"fff0117c", -- b690
		x"ff010001", -- b694
		x"3b7c0005", -- b698
		x"fffe4e4a", -- b69c
		x"4a6efffa", -- b6a0
		x"6600ff30", -- b6a4
		x"2b6f0008", -- b6a8
		x"fff6defc", -- b6ac
		x"000c4efa", -- b6b0
		x"00302c5f", -- b6b4
		x"2b5ffff6", -- b6b8
		x"70ffb06d", -- b6bc
		x"fffe6600", -- b6c0
		x"000a426e", -- b6c4
		x"000c6000", -- b6c8
		x"001870fe", -- b6cc
		x"b06dfffe", -- b6d0
		x"6600000c", -- b6d4
		x"3d7c0001", -- b6d8
		x"000c6000", -- b6dc
		x"00044e4a", -- b6e0
		x"4e5e2e9f", -- b6e4
		x"4e750000", -- b6e8
		x"4e56ffec", -- b6ec
		x"3d7c0003", -- b6f0
		x"001a2f2d", -- b6f4
		x"fff62f0e", -- b6f8
		x"487a01e8", -- b6fc
		x"2b4ffff6", -- b700
		x"2d6e0016", -- b704
		x"fff8206e", -- b708
		x"fff82d68", -- b70c
		x"0002fff4", -- b710
		x"226efff4", -- b714
		x"d3fc0000", -- b718
		x"800043d1", -- b71c
		x"2d49fff0", -- b720
		x"3d7c0001", -- b724
		x"fffe302e", -- b728
		x"fffe5340", -- b72c
		x"e340323b", -- b730
		x"00064efb", -- b734
		x"1002000a", -- b738
		x"003a0062", -- b73c
		x"00c00188", -- b740
		x"206efff4", -- b744
		x"08280006", -- b748
		x"000356c0", -- b74c
		x"44004a00", -- b750
		x"67000014", -- b754
		x"486effee", -- b758
		x"2f2e0016", -- b75c
		x"4ebaf8d6", -- b760
		x"3d6effee", -- b764
		x"fffc3d7c", -- b768
		x"0002fffe", -- b76c
		x"6000015e", -- b770
		x"558f2f2e", -- b774
		x"00162f2e", -- b778
		x"00084eba", -- b77c
		x"fc5a4a1f", -- b780
		x"6700000c", -- b784
		x"3d7c0004", -- b788
		x"fffe6000", -- b78c
		x"00083d7c", -- b790
		x"0003fffe", -- b794
		x"60000136", -- b798
		x"206efff4", -- b79c
		x"08280006", -- b7a0
		x"000356c0", -- b7a4
		x"44004a00", -- b7a8
		x"6700002e", -- b7ac
		x"486effee", -- b7b0
		x"2f2e0016", -- b7b4
		x"4ebaf87e", -- b7b8
		x"3d6effee", -- b7bc
		x"fffc082e", -- b7c0
		x"0002fffc", -- b7c4
		x"56c04400", -- b7c8
		x"4a006700", -- b7cc
		x"00083d7c", -- b7d0
		x"0002fffe", -- b7d4
		x"6000001c", -- b7d8
		x"558f2f2e", -- b7dc
		x"00124eba", -- b7e0
		x"9a744a1f", -- b7e4
		x"6700000c", -- b7e8
		x"3d7c0002", -- b7ec
		x"001a426e", -- b7f0
		x"fffe6000", -- b7f4
		x"00d8302e", -- b7f8
		x"0010907c", -- b7fc
		x"00816d00", -- b800
		x"00b4b07c", -- b804
		x"00016e00", -- b808
		x"00ace340", -- b80c
		x"323b0006", -- b810
		x"4efb1002", -- b814
		x"0004003a", -- b818
		x"206e0008", -- b81c
		x"2d50ffec", -- b820
		x"206effec", -- b824
		x"70001010", -- b828
		x"0c400081", -- b82c
		x"57c07202", -- b830
		x"b2680008", -- b834
		x"5fc1c200", -- b838
		x"6700000a", -- b83c
		x"426efffe", -- b840
		x"60000008", -- b844
		x"3d7c0005", -- b848
		x"fffe6000", -- b84c
		x"006e206e", -- b850
		x"00082d50", -- b854
		x"ffec206e", -- b858
		x"fff843e8", -- b85c
		x"000e2479", -- b860
		x"fffffed4", -- b864
		x"7206b30a", -- b868
		x"6600000a", -- b86c
		x"538166f6", -- b870
		x"70016002", -- b874
		x"4280226e", -- b878
		x"ffec7200", -- b87c
		x"12110c41", -- b880
		x"008257c1", -- b884
		x"c2002029", -- b888
		x"0002b0ae", -- b88c
		x"000c57c0", -- b890
		x"c0013229", -- b894
		x"0006b268", -- b898
		x"001457c1", -- b89c
		x"c2006700", -- b8a0
		x"000a426e", -- b8a4
		x"fffe6000", -- b8a8
		x"00083d7c", -- b8ac
		x"0005fffe", -- b8b0
		x"60000008", -- b8b4
		x"3d7c0005", -- b8b8
		x"fffe6000", -- b8bc
		x"00102f2e", -- b8c0
		x"00164eba", -- b8c4
		x"fa943d7c", -- b8c8
		x"0001fffe", -- b8cc
		x"4a6efffe", -- b8d0
		x"6600fe54", -- b8d4
		x"2b6f0008", -- b8d8
		x"fff6defc", -- b8dc
		x"000c4efa", -- b8e0
		x"001c2c5f", -- b8e4
		x"2b5ffff6", -- b8e8
		x"70ffb06d", -- b8ec
		x"fffe6600", -- b8f0
		x"000a426e", -- b8f4
		x"001a6000", -- b8f8
		x"00044e4a", -- b8fc
		x"4e5e205f", -- b900
		x"defc0012", -- b904
		x"4ed00000", -- b908
		x"4e56fff8", -- b90c
		x"422e0008", -- b910
		x"2d79ffff", -- b914
		x"fed4fff8", -- b918
		x"206efff8", -- b91c
		x"2d680010", -- b920
		x"fffc06ae", -- b924
		x"00000012", -- b928
		x"fffc558f", -- b92c
		x"2f2efffc", -- b930
		x"70001028", -- b934
		x"00603f00", -- b938
		x"4ebaf5b8", -- b93c
		x"1d5f0008", -- b940
		x"4e5e4e75", -- b944
		x"00004e56", -- b948
		x"fffc206e", -- b94c
		x"000830bc", -- b950
		x"00087001", -- b954
		x"b06e0014", -- b958
		x"66000026", -- b95c
		x"206e000c", -- b960
		x"2d50fffc", -- b964
		x"206efffc", -- b968
		x"10bcff03", -- b96c
		x"117cff00", -- b970
		x"000142a8", -- b974
		x"0002226e", -- b978
		x"00103169", -- b97c
		x"00140006", -- b980
		x"4e5e205f", -- b984
		x"defc000e", -- b988
		x"4ed00000", -- b98c
		x"4e56fffc", -- b990
		x"206e0008", -- b994
		x"30bc000a", -- b998
		x"7001b06e", -- b99c
		x"001a6600", -- b9a0
		x"002e206e", -- b9a4
		x"00122d50", -- b9a8
		x"fffc206e", -- b9ac
		x"fffc10bc", -- b9b0
		x"ff02117c", -- b9b4
		x"ff000001", -- b9b8
		x"216e000e", -- b9bc
		x"0002226e", -- b9c0
		x"00163169", -- b9c4
		x"00140006", -- b9c8
		x"316e000c", -- b9cc
		x"00084e5e", -- b9d0
		x"205fdefc", -- b9d4
		x"00144ed0", -- b9d8
		x"00004e56", -- b9dc
		x"fff4206e", -- b9e0
		x"000c7000", -- b9e4
		x"1010721e", -- b9e8
		x"d2405241", -- b9ec
		x"206e0008", -- b9f0
		x"3081206e", -- b9f4
		x"000c4a10", -- b9f8
		x"66000008", -- b9fc
		x"206e0008", -- ba00
		x"53507001", -- ba04
		x"b06e0018", -- ba08
		x"6600005a", -- ba0c
		x"206e0010", -- ba10
		x"2d50fff8", -- ba14
		x"2d79ffff", -- ba18
		x"fed4fff4", -- ba1c
		x"206efff8", -- ba20
		x"10bcff01", -- ba24
		x"117cff00", -- ba28
		x"0001226e", -- ba2c
		x"00142169", -- ba30
		x"00160002", -- ba34
		x"226e0014", -- ba38
		x"31690014", -- ba3c
		x"0006317c", -- ba40
		x"00020008", -- ba44
		x"4cba1e3f", -- ba48
		x"002648a8", -- ba4c
		x"1e3f000a", -- ba50
		x"226e000c", -- ba54
		x"45d1101a", -- ba58
		x"43e8001e", -- ba5c
		x"12c012da", -- ba60
		x"530062fa", -- ba64
		x"4e5e205f", -- ba68
		x"defc0012", -- ba6c
		x"4ed04850", -- ba70
		x"53333030", -- ba74
		x"20202020", -- ba78
		x"20202020", -- ba7c
		x"20202020", -- ba80
		x"20200000", -- ba84
		x"4e56fff0", -- ba88
		x"4a6e0018", -- ba8c
		x"66000028", -- ba90
		x"206e000c", -- ba94
		x"7018d050", -- ba98
		x"206e0008", -- ba9c
		x"3080206e", -- baa0
		x"0008703c", -- baa4
		x"b0506f00", -- baa8
		x"000a206e", -- baac
		x"000830bc", -- bab0
		x"003c6000", -- bab4
		x"00c87001", -- bab8
		x"b06e0018", -- babc
		x"660000be", -- bac0
		x"2d6e0014", -- bac4
		x"fff8206e", -- bac8
		x"fff82268", -- bacc
		x"0002d3fc", -- bad0
		x"00008000", -- bad4
		x"43d12d49", -- bad8
		x"fff4226e", -- badc
		x"fff445e9", -- bae0
		x"3ce02d4a", -- bae4
		x"fffc246e", -- bae8
		x"000c7018", -- baec
		x"d052246e", -- baf0
		x"00083480", -- baf4
		x"2d6efffc", -- baf8
		x"fff0246e", -- bafc
		x"fff02679", -- bb00
		x"fffffed4", -- bb04
		x"4c931300", -- bb08
		x"48921300", -- bb0c
		x"206efff8", -- bb10
		x"4ca81a00", -- bb14
		x"000848aa", -- bb18
		x"1a000006", -- bb1c
		x"226e0008", -- bb20
		x"700e9051", -- bb24
		x"44403540", -- bb28
		x"000c157c", -- bb2c
		x"00f8000e", -- bb30
		x"157c00f8", -- bb34
		x"000f157c", -- bb38
		x"00030010", -- bb3c
		x"157c0000", -- bb40
		x"0011157c", -- bb44
		x"00000012", -- bb48
		x"157c0000", -- bb4c
		x"0013357c", -- bb50
		x"06080014", -- bb54
		x"357c0609", -- bb58
		x"0016226e", -- bb5c
		x"001022ae", -- bb60
		x"fffc0691", -- bb64
		x"00000018", -- bb68
		x"226e0008", -- bb6c
		x"703cb051", -- bb70
		x"6f00000a", -- bb74
		x"226e0008", -- bb78
		x"32bc003c", -- bb7c
		x"4e5e205f", -- bb80
		x"defc0012", -- bb84
		x"4ed00001", -- bb88
		x"4e56fffc", -- bb8c
		x"0c798000", -- bb90
		x"fffffdd2", -- bb94
		x"57c00c79", -- bb98
		x"1000ffff", -- bb9c
		x"fdde57c1", -- bba0
		x"c2004a79", -- bba4
		x"fffffde0", -- bba8
		x"57c0c001", -- bbac
		x"4a79ffff", -- bbb0
		x"fde857c1", -- bbb4
		x"c2007001", -- bbb8
		x"b0b9ffff", -- bbbc
		x"fde25fc0", -- bbc0
		x"c0017201", -- bbc4
		x"b2b9ffff", -- bbc8
		x"fdda57c1", -- bbcc
		x"7402b4b9", -- bbd0
		x"fffffdda", -- bbd4
		x"57c28401", -- bbd8
		x"c4006700", -- bbdc
		x"002c1d7c", -- bbe0
		x"0001000c", -- bbe4
		x"2d79ffff", -- bbe8
		x"fed4fffc", -- bbec
		x"206efffc", -- bbf0
		x"2179ffff", -- bbf4
		x"fdda0062", -- bbf8
		x"2179ffff", -- bbfc
		x"fde20066", -- bc00
		x"42a8006a", -- bc04
		x"60000006", -- bc08
		x"422e000c", -- bc0c
		x"4e5e2e9f", -- bc10
		x"4e750001", -- bc14
		x"4e56fff0", -- bc18
		x"422efff9", -- bc1c
		x"2d79ffff", -- bc20
		x"fed4fff4", -- bc24
		x"206efff4", -- bc28
		x"3d680064", -- bc2c
		x"fffa2028", -- bc30
		x"0062d0a8", -- bc34
		x"00663d40", -- bc38
		x"fffc302e", -- bc3c
		x"fffa48c0", -- bc40
		x"2f002f3c", -- bc44
		x"00000100", -- bc48
		x"4879ffff", -- bc4c
		x"fdd21f3c", -- bc50
		x"ff014eba", -- bc54
		x"0888426e", -- bc58
		x"fffe302e", -- bc5c
		x"fffe48c0", -- bc60
		x"eb8041f9", -- bc64
		x"fffffdd2", -- bc68
		x"41f00800", -- bc6c
		x"2d48fff0", -- bc70
		x"206efff0", -- bc74
		x"70ffb068", -- bc78
		x"000a6600", -- bc7c
		x"000c3d7c", -- bc80
		x"0063fffe", -- bc84
		x"60000114", -- bc88
		x"206efff0", -- bc8c
		x"4a68000a", -- bc90
		x"6600000a", -- bc94
		x"526efffe", -- bc98
		x"60000100", -- bc9c
		x"4a2efff9", -- bca0
		x"6700007c", -- bca4
		x"206efff0", -- bca8
		x"3028001a", -- bcac
		x"02800000", -- bcb0
		x"7fff7201", -- bcb4
		x"b28057c0", -- bcb8
		x"08280007", -- bcbc
		x"001a56c1", -- bcc0
		x"4401c001", -- bcc4
		x"226e0008", -- bcc8
		x"24690008", -- bccc
		x"3212b268", -- bcd0
		x"000a57c1", -- bcd4
		x"c200246e", -- bcd8
		x"fff4202a", -- bcdc
		x"006eb0a8", -- bce0
		x"000c57c0", -- bce4
		x"c0012228", -- bce8
		x"0010e181", -- bcec
		x"2669000c", -- bcf0
		x"b29357c1", -- bcf4
		x"c2002669", -- bcf8
		x"00102013", -- bcfc
		x"b0a8001c", -- bd00
		x"57c0c001", -- bd04
		x"6700000a", -- bd08
		x"526efffe", -- bd0c
		x"6000000c", -- bd10
		x"3d7c0063", -- bd14
		x"fffe422e", -- bd18
		x"fff96000", -- bd1c
		x"007e206e", -- bd20
		x"00082268", -- bd24
		x"000870ff", -- bd28
		x"b05157c0", -- bd2c
		x"226efff0", -- bd30
		x"24680008", -- bd34
		x"3212b269", -- bd38
		x"000a57c1", -- bd3c
		x"82003029", -- bd40
		x"001a0280", -- bd44
		x"00007fff", -- bd48
		x"7401b480", -- bd4c
		x"57c00829", -- bd50
		x"0007001a", -- bd54
		x"56c24402", -- bd58
		x"c002c200", -- bd5c
		x"67000036", -- bd60
		x"24680008", -- bd64
		x"34a9000a", -- bd68
		x"246efff4", -- bd6c
		x"2569000c", -- bd70
		x"006e2029", -- bd74
		x"0010e180", -- bd78
		x"2668000c", -- bd7c
		x"26802668", -- bd80
		x"001026a9", -- bd84
		x"001c1d7c", -- bd88
		x"0001fff9", -- bd8c
		x"526efffe", -- bd90
		x"60000008", -- bd94
		x"3d7c0063", -- bd98
		x"fffe7007", -- bd9c
		x"b06efffe", -- bda0
		x"6c00feb8", -- bda4
		x"7063b06e", -- bda8
		x"fffe6600", -- bdac
		x"000c3d6e", -- bdb0
		x"fffcfffa", -- bdb4
		x"60000006", -- bdb8
		x"526efffa", -- bdbc
		x"302efffa", -- bdc0
		x"b06efffc", -- bdc4
		x"6d00fe74", -- bdc8
		x"1d6efff9", -- bdcc
		x"000c4e5e", -- bdd0
		x"2e9f4e75", -- bdd4
		x"00004e56", -- bdd8
		x"ffda422e", -- bddc
		x"00182079", -- bde0
		x"fffffed4", -- bde4
		x"2d680010", -- bde8
		x"fffc06ae", -- bdec
		x"00000012", -- bdf0
		x"fffc2d79", -- bdf4
		x"fffffed4", -- bdf8
		x"ffe22d6e", -- bdfc
		x"fffcffde", -- be00
		x"558f2f2e", -- be04
		x"fffc206e", -- be08
		x"ffe27000", -- be0c
		x"10280060", -- be10
		x"3f004eba", -- be14
		x"f0de4a1f", -- be18
		x"6600000a", -- be1c
		x"3b7c0003", -- be20
		x"fffe4e4a", -- be24
		x"206e0014", -- be28
		x"43fa03ac", -- be2c
		x"70001010", -- be30
		x"5240b109", -- be34
		x"6600000e", -- be38
		x"534066f6", -- be3c
		x"3b7c0003", -- be40
		x"fffe4e4a", -- be44
		x"206effe2", -- be48
		x"217cffff", -- be4c
		x"ffff006e", -- be50
		x"226effde", -- be54
		x"7000246e", -- be58
		x"00141012", -- be5c
		x"23400016", -- be60
		x"48690016", -- be64
		x"4eba93b4", -- be68
		x"206effde", -- be6c
		x"42680014", -- be70
		x"42672f2e", -- be74
		x"fffc486e", -- be78
		x"fff42f2e", -- be7c
		x"0014486e", -- be80
		x"fffa4eba", -- be84
		x"fb564267", -- be88
		x"2f2efffc", -- be8c
		x"486efff4", -- be90
		x"486efffa", -- be94
		x"486efff8", -- be98
		x"4ebafbea", -- be9c
		x"3d7c0001", -- bea0
		x"ffee3d7c", -- bea4
		x"0008fff2", -- bea8
		x"2d7c0000", -- beac
		x"0006ffe6", -- beb0
		x"302effee", -- beb4
		x"5340e340", -- beb8
		x"323b0006", -- bebc
		x"4efb1002", -- bec0
		x"000600a6", -- bec4
		x"016e2f2e", -- bec8
		x"fffc3f2e", -- becc
		x"fff84eba", -- bed0
		x"f0ca3f3c", -- bed4
		x"00012f2e", -- bed8
		x"fffc486e", -- bedc
		x"fff4486e", -- bee0
		x"fffa486e", -- bee4
		x"fff84eba", -- bee8
		x"fb9c3f3c", -- beec
		x"00012f2e", -- bef0
		x"fffc486e", -- bef4
		x"fff42f2e", -- bef8
		x"0014486e", -- befc
		x"fffa4eba", -- bf00
		x"fada558f", -- bf04
		x"2f2efffc", -- bf08
		x"4ebaf666", -- bf0c
		x"3d5ffff0", -- bf10
		x"7003b06e", -- bf14
		x"fff057c0", -- bf18
		x"7204b26e", -- bf1c
		x"fff057c1", -- bf20
		x"82006700", -- bf24
		x"000c3d7c", -- bf28
		x"0002ffee", -- bf2c
		x"6000001a", -- bf30
		x"558f486e", -- bf34
		x"fff24eba", -- bf38
		x"182a4a1f", -- bf3c
		x"6600000a", -- bf40
		x"3b7c0005", -- bf44
		x"fffe4e4a", -- bf48
		x"2f3c000f", -- bf4c
		x"42402f2e", -- bf50
		x"ffe64eba", -- bf54
		x"c2582d5f", -- bf58
		x"ffea486e", -- bf5c
		x"ffea4eba", -- bf60
		x"92ba6000", -- bf64
		x"01e8558f", -- bf68
		x"2f2efffc", -- bf6c
		x"486effea", -- bf70
		x"3f3c0081", -- bf74
		x"2f3c0000", -- bf78
		x"0063486e", -- bf7c
		x"fff44eba", -- bf80
		x"f768301f", -- bf84
		x"e340323b", -- bf88
		x"00064efb", -- bf8c
		x"10020076", -- bf90
		x"009c0012", -- bf94
		x"00083d7c", -- bf98
		x"0003ffee", -- bf9c
		x"6000008c", -- bfa0
		x"558f486e", -- bfa4
		x"fff24eba", -- bfa8
		x"17ba4a1f", -- bfac
		x"6700000c", -- bfb0
		x"3d7c0001", -- bfb4
		x"ffee6000", -- bfb8
		x"0048206e", -- bfbc
		x"ffe20828", -- bfc0
		x"0002000a", -- bfc4
		x"56c04400", -- bfc8
		x"4a006700", -- bfcc
		x"002c3d7c", -- bfd0
		x"7ffffff2", -- bfd4
		x"226effde", -- bfd8
		x"1029000d", -- bfdc
		x"02000007", -- bfe0
		x"72001200", -- bfe4
		x"700ad240", -- bfe8
		x"48c12d41", -- bfec
		x"ffe63d7c", -- bff0
		x"0001ffee", -- bff4
		x"6000000a", -- bff8
		x"3b7c0002", -- bffc
		x"fffe4e4a", -- c000
		x"60000028", -- c004
		x"558f486e", -- c008
		x"fff24eba", -- c00c
		x"17564a1f", -- c010
		x"6700000c", -- c014
		x"3d7c0001", -- c018
		x"ffee6000", -- c01c
		x"000a3b7c", -- c020
		x"0004fffe", -- c024
		x"4e4a6000", -- c028
		x"00026000", -- c02c
		x"0120426e", -- c030
		x"ffee206e", -- c034
		x"ffde43e8", -- c038
		x"000e246e", -- c03c
		x"ffe27006", -- c040
		x"b30a6600", -- c044
		x"000a5380", -- c048
		x"66f66000", -- c04c
		x"000c3d7c", -- c050
		x"0002ffee", -- c054
		x"600000ee", -- c058
		x"2d6efff4", -- c05c
		x"ffda206e", -- c060
		x"ffda226e", -- c064
		x"ffde2029", -- c068
		x"0016b0a8", -- c06c
		x"00026700", -- c070
		x"000c3d7c", -- c074
		x"0002ffee", -- c078
		x"600000ca", -- c07c
		x"206effda", -- c080
		x"4a280001", -- c084
		x"66000056", -- c088
		x"226effde", -- c08c
		x"700ab069", -- c090
		x"001e6600", -- c094
		x"000c3d7c", -- c098
		x"0002ffee", -- c09c
		x"6000003a", -- c0a0
		x"206effda", -- c0a4
		x"43e8000a", -- c0a8
		x"246e0014", -- c0ac
		x"70001011", -- c0b0
		x"5240b30a", -- c0b4
		x"6600000a", -- c0b8
		x"534066f6", -- c0bc
		x"6000000c", -- c0c0
		x"3d7c0002", -- c0c4
		x"ffee6000", -- c0c8
		x"0010206e", -- c0cc
		x"ffda226e", -- c0d0
		x"ffde3368", -- c0d4
		x"00060014", -- c0d8
		x"6000006a", -- c0dc
		x"42aefff4", -- c0e0
		x"3d7c0002", -- c0e4
		x"ffee206e", -- c0e8
		x"ffda7004", -- c0ec
		x"b0280001", -- c0f0
		x"57c07205", -- c0f4
		x"b2280001", -- c0f8
		x"57c18200", -- c0fc
		x"67000034", -- c100
		x"526efff2", -- c104
		x"701090ae", -- c108
		x"ffe66c02", -- c10c
		x"5280e280", -- c110
		x"d1aeffe6", -- c114
		x"2f3c000f", -- c118
		x"42402f2e", -- c11c
		x"ffe64eba", -- c120
		x"c08c2d5f", -- c124
		x"ffea486e", -- c128
		x"ffea4eba", -- c12c
		x"90ee6000", -- c130
		x"0014206e", -- c134
		x"ffda701b", -- c138
		x"b0280001", -- c13c
		x"67000006", -- c140
		x"426effee", -- c144
		x"2f2efffc", -- c148
		x"4ebaf20e", -- c14c
		x"4a6effee", -- c150
		x"6600fd5e", -- c154
		x"4aaefff4", -- c158
		x"67000072", -- c15c
		x"206effe2", -- c160
		x"42a8006e", -- c164
		x"42a72f3c", -- c168
		x"00000100", -- c16c
		x"4879ffff", -- c170
		x"fdd21f3c", -- c174
		x"ff014eba", -- c178
		x"0364558f", -- c17c
		x"2f0e4eba", -- c180
		x"fa084a1f", -- c184
		x"6600003a", -- c188
		x"206e0008", -- c18c
		x"70ffb050", -- c190
		x"57c00200", -- c194
		x"00011d40", -- c198
		x"0018206e", -- c19c
		x"ffe242a8", -- c1a0
		x"006242a8", -- c1a4
		x"006e226e", -- c1a8
		x"00104291", -- c1ac
		x"226e000c", -- c1b0
		x"22bcffff", -- c1b4
		x"ffff226e", -- c1b8
		x"00084251", -- c1bc
		x"6000000e", -- c1c0
		x"558f2f0e", -- c1c4
		x"4ebafa4e", -- c1c8
		x"1d5f0018", -- c1cc
		x"4e5e205f", -- c1d0
		x"defc0010", -- c1d4
		x"4ed00000", -- c1d8
		x"00014e56", -- c1dc
		x"fffc206e", -- c1e0
		x"00083028", -- c1e4
		x"fff20240", -- c1e8
		x"000f5240", -- c1ec
		x"3140fff2", -- c1f0
		x"22680008", -- c1f4
		x"2469fff0", -- c1f8
		x"246a0002", -- c1fc
		x"3028fff2", -- c200
		x"48c0e780", -- c204
		x"d5fc0000", -- c208
		x"801045f2", -- c20c
		x"08002d4a", -- c210
		x"fffc42a8", -- c214
		x"ffea246e", -- c218
		x"fffc3012", -- c21c
		x"3140ffec", -- c220
		x"116a0003", -- c224
		x"ffeb4e5e", -- c228
		x"2e9f4e75", -- c22c
		x"00014e56", -- c230
		x"ffe2206e", -- c234
		x"00082d68", -- c238
		x"fff0ffe6", -- c23c
		x"3d7c0001", -- c240
		x"fff4302e", -- c244
		x"fff45340", -- c248
		x"e340323b", -- c24c
		x"00064efb", -- c250
		x"10020008", -- c254
		x"00500110", -- c258
		x"01664267", -- c25c
		x"206e0008", -- c260
		x"2f28fff0", -- c264
		x"4868ffec", -- c268
		x"2f28fff8", -- c26c
		x"3f2e000e", -- c270
		x"486efff8", -- c274
		x"4ebaf716", -- c278
		x"4267206e", -- c27c
		x"00082f28", -- c280
		x"fff04868", -- c284
		x"ffec486e", -- c288
		x"fff8486e", -- c28c
		x"fffa4eba", -- c290
		x"f7f43d7c", -- c294
		x"000afff6", -- c298
		x"3d7c0002", -- c29c
		x"fff46000", -- c2a0
		x"022a206e", -- c2a4
		x"00082f28", -- c2a8
		x"fff03f2e", -- c2ac
		x"fffa4eba", -- c2b0
		x"ecea3f3c", -- c2b4
		x"0001206e", -- c2b8
		x"00082f28", -- c2bc
		x"fff04868", -- c2c0
		x"ffec486e", -- c2c4
		x"fff8486e", -- c2c8
		x"fffa4eba", -- c2cc
		x"f7b83f3c", -- c2d0
		x"0001206e", -- c2d4
		x"00082f28", -- c2d8
		x"fff04868", -- c2dc
		x"ffec2f28", -- c2e0
		x"fff83f2e", -- c2e4
		x"000e486e", -- c2e8
		x"fff84eba", -- c2ec
		x"f6a0558f", -- c2f0
		x"206e0008", -- c2f4
		x"2f28fff0", -- c2f8
		x"4ebaf276", -- c2fc
		x"301f48c0", -- c300
		x"2d40fffc", -- c304
		x"7003b0ae", -- c308
		x"fffc57c0", -- c30c
		x"7204b2ae", -- c310
		x"fffc57c1", -- c314
		x"82006700", -- c318
		x"000c3d7c", -- c31c
		x"0003fff4", -- c320
		x"6000001a", -- c324
		x"558f486e", -- c328
		x"fff64eba", -- c32c
		x"14364a1f", -- c330
		x"6600000a", -- c334
		x"3b7c0005", -- c338
		x"fffe4e4a", -- c33c
		x"2f3c000f", -- c340
		x"4240700a", -- c344
		x"906efff6", -- c348
		x"564048c0", -- c34c
		x"2f004eba", -- c350
		x"be5c2d5f", -- c354
		x"ffee486e", -- c358
		x"ffee4eba", -- c35c
		x"8ebe6000", -- c360
		x"016a558f", -- c364
		x"206e0008", -- c368
		x"2f28fff0", -- c36c
		x"486effee", -- c370
		x"3f3c0082", -- c374
		x"2f28fff8", -- c378
		x"4868ffec", -- c37c
		x"4ebaf36a", -- c380
		x"7003b05f", -- c384
		x"6600000c", -- c388
		x"3d7c0004", -- c38c
		x"fff46000", -- c390
		x"0024558f", -- c394
		x"486efff6", -- c398
		x"4eba13c8", -- c39c
		x"4a1f6700", -- c3a0
		x"000c3d7c", -- c3a4
		x"0002fff4", -- c3a8
		x"6000000a", -- c3ac
		x"3b7c0004", -- c3b0
		x"fffe4e4a", -- c3b4
		x"60000114", -- c3b8
		x"426efff4", -- c3bc
		x"206e0008", -- c3c0
		x"2d68ffec", -- c3c4
		x"ffe2226e", -- c3c8
		x"ffe245e9", -- c3cc
		x"00082d4a", -- c3d0
		x"ffea246e", -- c3d4
		x"ffe63d6a", -- c3d8
		x"0006fff2", -- c3dc
		x"516a001e", -- c3e0
		x"4a290001", -- c3e4
		x"57c0322a", -- c3e8
		x"001e48c1", -- c3ec
		x"b2ae000c", -- c3f0
		x"5fc1c200", -- c3f4
		x"6700009c", -- c3f8
		x"302a001e", -- c3fc
		x"48c091ae", -- c400
		x"000c4aae", -- c404
		x"000c6f00", -- c408
		x"00083d7c", -- c40c
		x"0001fff4", -- c410
		x"206effe6", -- c414
		x"51680020", -- c418
		x"206effe6", -- c41c
		x"4a68001e", -- c420
		x"6f00006c", -- c424
		x"2f2effea", -- c428
		x"226e0008", -- c42c
		x"2f29000a", -- c430
		x"30280020", -- c434
		x"48c02f00", -- c438
		x"4eba1310", -- c43c
		x"206effe6", -- c440
		x"30280020", -- c444
		x"9168001e", -- c448
		x"226e0008", -- c44c
		x"30280020", -- c450
		x"48c0d1a9", -- c454
		x"fff83028", -- c458
		x"002048c0", -- c45c
		x"d1a9000a", -- c460
		x"4a68001e", -- c464
		x"6f000026", -- c468
		x"0c6803c4", -- c46c
		x"001e6f00", -- c470
		x"000c317c", -- c474
		x"03c40020", -- c478
		x"6000000c", -- c47c
		x"206effe6", -- c480
		x"3168001e", -- c484
		x"00202f0e", -- c488
		x"4ebafd50", -- c48c
		x"608a6000", -- c490
		x"002e206e", -- c494
		x"ffe27002", -- c498
		x"b0280001", -- c49c
		x"57c07203", -- c4a0
		x"b2280001", -- c4a4
		x"57c18200", -- c4a8
		x"6700000e", -- c4ac
		x"3b7c0004", -- c4b0
		x"fffe4e4a", -- c4b4
		x"60000008", -- c4b8
		x"3d7c0003", -- c4bc
		x"fff4206e", -- c4c0
		x"00082f28", -- c4c4
		x"fff04eba", -- c4c8
		x"ee904a6e", -- c4cc
		x"fff46600", -- c4d0
		x"fd724e5e", -- c4d4
		x"205f504f", -- c4d8
		x"4ed00000", -- c4dc
		x"4e56ffec", -- c4e0
		x"2079ffff", -- c4e4
		x"fed44aa8", -- c4e8
		x"006e6c00", -- c4ec
		x"000a3b7c", -- c4f0
		x"0003fffe", -- c4f4
		x"4e4a2079", -- c4f8
		x"fffffed4", -- c4fc
		x"2d680010", -- c500
		x"fff006ae", -- c504
		x"00000012", -- c508
		x"fff02d7c", -- c50c
		x"000005ca", -- c510
		x"fffc4a2e", -- c514
		x"00086600", -- c518
		x"00102079", -- c51c
		x"fffffed4", -- c520
		x"2028006e", -- c524
		x"d1ae0012", -- c528
		x"202e0012", -- c52c
		x"e1802d40", -- c530
		x"fff84aae", -- c534
		x"000e6f00", -- c538
		x"0032202e", -- c53c
		x"000eb0ae", -- c540
		x"fffc6e00", -- c544
		x"000c2d6e", -- c548
		x"000efff4", -- c54c
		x"60000008", -- c550
		x"2d6efffc", -- c554
		x"fff42f2e", -- c558
		x"fff42f0e", -- c55c
		x"4ebafcd0", -- c560
		x"202efff4", -- c564
		x"91ae000e", -- c568
		x"60c84e5e", -- c56c
		x"205fdefc", -- c570
		x"000e4ed0", -- c574
		x"00004e56", -- c578
		x"ffec1d7c", -- c57c
		x"0001fff2", -- c580
		x"1d7c0001", -- c584
		x"fff32d6e", -- c588
		x"0008ffec", -- c58c
		x"42672f2e", -- c590
		x"0008486e", -- c594
		x"fff8486e", -- c598
		x"fffe4eba", -- c59c
		x"f3aa4267", -- c5a0
		x"2f2e0008", -- c5a4
		x"486efff8", -- c5a8
		x"486efffe", -- c5ac
		x"486efffc", -- c5b0
		x"4ebaf4d2", -- c5b4
		x"3d7c0003", -- c5b8
		x"fff42f2e", -- c5bc
		x"00083f2e", -- c5c0
		x"fffc4eba", -- c5c4
		x"e9d63f3c", -- c5c8
		x"00012f2e", -- c5cc
		x"0008486e", -- c5d0
		x"fff8486e", -- c5d4
		x"fffe486e", -- c5d8
		x"fffc4eba", -- c5dc
		x"f4a83f3c", -- c5e0
		x"00012f2e", -- c5e4
		x"0008486e", -- c5e8
		x"fff8486e", -- c5ec
		x"fffe4eba", -- c5f0
		x"f356558f", -- c5f4
		x"2f2e0008", -- c5f8
		x"4ebaef76", -- c5fc
		x"3d5ffff6", -- c600
		x"7003b06e", -- c604
		x"fff66600", -- c608
		x"000c1d7c", -- c60c
		x"0001fff1", -- c610
		x"60000038", -- c614
		x"558f486e", -- c618
		x"fff44eba", -- c61c
		x"11464a1f", -- c620
		x"6700001e", -- c624
		x"4a2efff3", -- c628
		x"67000012", -- c62c
		x"7001b06e", -- c630
		x"fff657c0", -- c634
		x"0200ff01", -- c638
		x"1d40fff3", -- c63c
		x"6000000c", -- c640
		x"422efff2", -- c644
		x"1d7cff01", -- c648
		x"fff14a2e", -- c64c
		x"fff16700", -- c650
		x"ff6a4a2e", -- c654
		x"fff26700", -- c658
		x"001e4a2e", -- c65c
		x"fff36700", -- c660
		x"000c3d7c", -- c664
		x"0003000c", -- c668
		x"60000008", -- c66c
		x"3d7c0004", -- c670
		x"000c6000", -- c674
		x"00184a2e", -- c678
		x"fff36700", -- c67c
		x"000c3d7c", -- c680
		x"0001000c", -- c684
		x"60000006", -- c688
		x"426e000c", -- c68c
		x"206effec", -- c690
		x"42680014", -- c694
		x"2279ffff", -- c698
		x"fed4237c", -- c69c
		x"ffffffff", -- c6a0
		x"006e4e5e", -- c6a4
		x"2e9f4e75", -- c6a8
		x"00004e56", -- c6ac
		x"fffa2079", -- c6b0
		x"fffffed4", -- c6b4
		x"2d680010", -- c6b8
		x"fffc06ae", -- c6bc
		x"00000012", -- c6c0
		x"fffc2f2d", -- c6c4
		x"fff62f0e", -- c6c8
		x"487a002e", -- c6cc
		x"2b4ffff6", -- c6d0
		x"206efffc", -- c6d4
		x"4a680014", -- c6d8
		x"6f000010", -- c6dc
		x"558f2f2e", -- c6e0
		x"fffc4eba", -- c6e4
		x"fe923d5f", -- c6e8
		x"fffa2b6f", -- c6ec
		x"0008fff6", -- c6f0
		x"defc000c", -- c6f4
		x"4efa0008", -- c6f8
		x"2c5f2b5f", -- c6fc
		x"fff64e5e", -- c700
		x"4e750000", -- c704
		x"4e56fff2", -- c708
		x"2d79ffff", -- c70c
		x"fed4fffa", -- c710
		x"2d6e0008", -- c714
		x"fff6206e", -- c718
		x"fffa226e", -- c71c
		x"fff62368", -- c720
		x"0336001a", -- c724
		x"422effff", -- c728
		x"206efff6", -- c72c
		x"4aa8001a", -- c730
		x"56c0122e", -- c734
		x"ffff0841", -- c738
		x"0000c001", -- c73c
		x"67000030", -- c740
		x"226efffa", -- c744
		x"2468001a", -- c748
		x"70001029", -- c74c
		x"0060b052", -- c750
		x"6600000c", -- c754
		x"1d7c0001", -- c758
		x"ffff6000", -- c75c
		x"0010206e", -- c760
		x"fff62268", -- c764
		x"001a2169", -- c768
		x"0004001a", -- c76c
		x"60ba4a2e", -- c770
		x"ffff6600", -- c774
		x"003e206e", -- c778
		x"fff64868", -- c77c
		x"001a2f3c", -- c780
		x"00000188", -- c784
		x"4eba0fb2", -- c788
		x"206efff6", -- c78c
		x"2d68001a", -- c790
		x"fff2226e", -- c794
		x"fffa246e", -- c798
		x"fff27000", -- c79c
		x"10290060", -- c7a0
		x"3480426a", -- c7a4
		x"00022569", -- c7a8
		x"03360004", -- c7ac
		x"2368001a", -- c7b0
		x"03364e5e", -- c7b4
		x"2e9f4e75", -- c7b8
		x"00004e56", -- c7bc
		x"fff42d79", -- c7c0
		x"fffffed4", -- c7c4
		x"fff8206e", -- c7c8
		x"fff82d68", -- c7cc
		x"0010fffc", -- c7d0
		x"06ae0000", -- c7d4
		x"0012fffc", -- c7d8
		x"226e000a", -- c7dc
		x"42114a2e", -- c7e0
		x"00126700", -- c7e4
		x"003a217a", -- c7e8
		x"e2ce005e", -- c7ec
		x"226e000e", -- c7f0
		x"22a8005e", -- c7f4
		x"558f2f2e", -- c7f8
		x"fffc7000", -- c7fc
		x"10280060", -- c800
		x"3f004eba", -- c804
		x"e6ee206e", -- c808
		x"000a109f", -- c80c
		x"206e000a", -- c810
		x"4a106700", -- c814
		x"000a2f2e", -- c818
		x"fffc4eba", -- c81c
		x"fee82d6e", -- c820
		x"fffcfff4", -- c824
		x"206efff4", -- c828
		x"216e000e", -- c82c
		x"0022317c", -- c830
		x"00010026", -- c834
		x"226efff8", -- c838
		x"137cff03", -- c83c
		x"0061206e", -- c840
		x"000a1d50", -- c844
		x"00164e5e", -- c848
		x"205fdefc", -- c84c
		x"000e4ed0", -- c850
		x"00004e56", -- c854
		x"fff0206e", -- c858
		x"000a4210", -- c85c
		x"2d79ffff", -- c860
		x"fed4fff8", -- c864
		x"206efff8", -- c868
		x"43e8005e", -- c86c
		x"2d49fff4", -- c870
		x"2d680010", -- c874
		x"fffc06ae", -- c878
		x"00000012", -- c87c
		x"fffc226e", -- c880
		x"000a4211", -- c884
		x"4a2e0012", -- c888
		x"6700000c", -- c88c
		x"217ae224", -- c890
		x"005e6000", -- c894
		x"0018206e", -- c898
		x"fff47000", -- c89c
		x"10280002", -- c8a0
		x"52401140", -- c8a4
		x"0002117c", -- c8a8
		x"00000001", -- c8ac
		x"206efff4", -- c8b0
		x"7020b028", -- c8b4
		x"000252c0", -- c8b8
		x"226e000a", -- c8bc
		x"12110841", -- c8c0
		x"0000c200", -- c8c4
		x"67000042", -- c8c8
		x"558f2f2e", -- c8cc
		x"fffc7000", -- c8d0
		x"10280002", -- c8d4
		x"3f004eba", -- c8d8
		x"e61a206e", -- c8dc
		x"000a109f", -- c8e0
		x"206e000a", -- c8e4
		x"4a106700", -- c8e8
		x"000e2f2e", -- c8ec
		x"fffc4eba", -- c8f0
		x"fe146000", -- c8f4
		x"0012206e", -- c8f8
		x"fff47000", -- c8fc
		x"10280002", -- c900
		x"52401140", -- c904
		x"000260a4", -- c908
		x"206efff8", -- c90c
		x"226e000e", -- c910
		x"22a8005e", -- c914
		x"2d6efffc", -- c918
		x"fff0226e", -- c91c
		x"fff0236e", -- c920
		x"000e0022", -- c924
		x"337c0001", -- c928
		x"0026117c", -- c92c
		x"00030061", -- c930
		x"206e000a", -- c934
		x"1d500016", -- c938
		x"4e5e205f", -- c93c
		x"defc000e", -- c940
		x"4ed00100", -- c944
		x"02120203", -- c948
		x"01010304", -- c94c
		x"16020405", -- c950
		x"15050503", -- c954
		x"06060607", -- c958
		x"02000708", -- c95c
		x"0f100809", -- c960
		x"070e030a", -- c964
		x"0b080408", -- c968
		x"1408090c", -- c96c
		x"0d080a00", -- c970
		x"00000b06", -- c974
		x"11080107", -- c978
		x"0e070108", -- c97c
		x"0e070106", -- c980
		x"10060c06", -- c984
		x"00000d01", -- c988
		x"00000e08", -- c98c
		x"04000f0c", -- c990
		x"130e0f0c", -- c994
		x"05011002", -- c998
		x"00000001", -- c99c
		x"4e56fff6", -- c9a0
		x"1d7c0001", -- c9a4
		x"ffff206e", -- c9a8
		x"00082d68", -- c9ac
		x"fffcfff8", -- c9b0
		x"70013d68", -- c9b4
		x"ffeafff6", -- c9b8
		x"b06efff6", -- c9bc
		x"6e00003e", -- c9c0
		x"3d40fffc", -- c9c4
		x"206e0008", -- c9c8
		x"2268ffec", -- c9cc
		x"302efffc", -- c9d0
		x"c1fc0018", -- c9d4
		x"43f108e8", -- c9d8
		x"246efff8", -- c9dc
		x"47ea000e", -- c9e0
		x"7006b30b", -- c9e4
		x"6600000e", -- c9e8
		x"538066f6", -- c9ec
		x"422effff", -- c9f0
		x"6000000a", -- c9f4
		x"302efffc", -- c9f8
		x"524068bc", -- c9fc
		x"206e0008", -- ca00
		x"7010b068", -- ca04
		x"ffea5ec0", -- ca08
		x"c02effff", -- ca0c
		x"0200ff01", -- ca10
		x"1d40000c", -- ca14
		x"4e5e2e9f", -- ca18
		x"4e750001", -- ca1c
		x"4e56fff4", -- ca20
		x"2d79ffff", -- ca24
		x"fed4fff4", -- ca28
		x"4267206e", -- ca2c
		x"00082f28", -- ca30
		x"fffc4868", -- ca34
		x"fff42f28", -- ca38
		x"00084868", -- ca3c
		x"fffa4eba", -- ca40
		x"ef9a4267", -- ca44
		x"206e0008", -- ca48
		x"2f28fffc", -- ca4c
		x"4868fff4", -- ca50
		x"4868fffa", -- ca54
		x"4868fff8", -- ca58
		x"4ebaf02a", -- ca5c
		x"3d7c0002", -- ca60
		x"fffc1d7c", -- ca64
		x"0001fffa", -- ca68
		x"1d7c0001", -- ca6c
		x"fffb206e", -- ca70
		x"00082f28", -- ca74
		x"fffc3f28", -- ca78
		x"fff84eba", -- ca7c
		x"e51e3f3c", -- ca80
		x"0001206e", -- ca84
		x"00082f28", -- ca88
		x"fffc4868", -- ca8c
		x"fff44868", -- ca90
		x"fffa4868", -- ca94
		x"fff84eba", -- ca98
		x"efec3f3c", -- ca9c
		x"0001206e", -- caa0
		x"00082f28", -- caa4
		x"fffc4868", -- caa8
		x"fff42f28", -- caac
		x"00084868", -- cab0
		x"fffa4eba", -- cab4
		x"ef26558f", -- cab8
		x"206e0008", -- cabc
		x"2f28fffc", -- cac0
		x"4ebaeaae", -- cac4
		x"3d5ffffe", -- cac8
		x"7003b06e", -- cacc
		x"fffe6600", -- cad0
		x"000c1d7c", -- cad4
		x"0001fff9", -- cad8
		x"60000038", -- cadc
		x"558f486e", -- cae0
		x"fffc4eba", -- cae4
		x"0c7e4a1f", -- cae8
		x"6700001e", -- caec
		x"4a2efffb", -- caf0
		x"67000012", -- caf4
		x"7001b06e", -- caf8
		x"fffe57c0", -- cafc
		x"0200ff01", -- cb00
		x"1d40fffb", -- cb04
		x"6000000c", -- cb08
		x"422efffa", -- cb0c
		x"1d7cff01", -- cb10
		x"fff94a2e", -- cb14
		x"fff96700", -- cb18
		x"ff564a2e", -- cb1c
		x"fffa6700", -- cb20
		x"001e4a2e", -- cb24
		x"fffb6700", -- cb28
		x"000c3d7c", -- cb2c
		x"0003000c", -- cb30
		x"60000008", -- cb34
		x"3d7c0004", -- cb38
		x"000c6000", -- cb3c
		x"00184a2e", -- cb40
		x"fffb6700", -- cb44
		x"000c3d7c", -- cb48
		x"0001000c", -- cb4c
		x"60000006", -- cb50
		x"426e000c", -- cb54
		x"4e5e2e9f", -- cb58
		x"4e750000", -- cb5c
		x"4e56ffc0", -- cb60
		x"2079ffff", -- cb64
		x"fed42d68", -- cb68
		x"0010fffc", -- cb6c
		x"06ae0000", -- cb70
		x"0012fffc", -- cb74
		x"2d79ffff", -- cb78
		x"fed4ffcc", -- cb7c
		x"2d6efffc", -- cb80
		x"ffc841fa", -- cb84
		x"09021018", -- cb88
		x"246e0008", -- cb8c
		x"43d212c0", -- cb90
		x"12d85300", -- cb94
		x"62fa206e", -- cb98
		x"ffc82268", -- cb9c
		x"001a3d69", -- cba0
		x"0002ffea", -- cba4
		x"2268001a", -- cba8
		x"43e90008", -- cbac
		x"2d49ffec", -- cbb0
		x"422effd9", -- cbb4
		x"3d7c0003", -- cbb8
		x"fff2226e", -- cbbc
		x"ffcc7000", -- cbc0
		x"10290061", -- cbc4
		x"3d40ffe2", -- cbc8
		x"3d680026", -- cbcc
		x"fff01d7c", -- cbd0
		x"0001000c", -- cbd4
		x"2f2dfff6", -- cbd8
		x"2f0e487a", -- cbdc
		x"08742b4f", -- cbe0
		x"fff6302e", -- cbe4
		x"fff048c0", -- cbe8
		x"e58041fa", -- cbec
		x"fd56d0fc", -- cbf0
		x"fffd7200", -- cbf4
		x"12300800", -- cbf8
		x"3d41ffd0", -- cbfc
		x"302efff0", -- cc00
		x"48c0e580", -- cc04
		x"41fafd3c", -- cc08
		x"d0fcfffe", -- cc0c
		x"72001230", -- cc10
		x"08003d41", -- cc14
		x"ffd2302e", -- cc18
		x"fff048c0", -- cc1c
		x"e58041fa", -- cc20
		x"fd22d0fc", -- cc24
		x"ffff7200", -- cc28
		x"12300800", -- cc2c
		x"3d41ffd4", -- cc30
		x"302efff0", -- cc34
		x"48c0e580", -- cc38
		x"41fafd08", -- cc3c
		x"d0fcfffc", -- cc40
		x"72001230", -- cc44
		x"08005341", -- cc48
		x"6d0007d0", -- cc4c
		x"b27c000f", -- cc50
		x"6e0007c8", -- cc54
		x"e341303b", -- cc58
		x"10064efb", -- cc5c
		x"00020020", -- cc60
		x"00ca0126", -- cc64
		x"017e02d0", -- cc68
		x"03440396", -- cc6c
		x"046404c8", -- cc70
		x"055e065c", -- cc74
		x"06d40748", -- cc78
		x"07680790", -- cc7c
		x"07aa558f", -- cc80
		x"486effe2", -- cc84
		x"4eba0adc", -- cc88
		x"4a1f6700", -- cc8c
		x"0092206e", -- cc90
		x"ffcc4cba", -- cc94
		x"0e0007f2", -- cc98
		x"48900e00", -- cc9c
		x"43fa07e8", -- cca0
		x"101945e8", -- cca4
		x"00ce14c0", -- cca8
		x"14d95300", -- ccac
		x"62fa226e", -- ccb0
		x"ffc842a9", -- ccb4
		x"0016337c", -- ccb8
		x"ffff0014", -- ccbc
		x"302efff0", -- ccc0
		x"52403340", -- ccc4
		x"0026558f", -- ccc8
		x"2f0e4eba", -- cccc
		x"fd50301f", -- ccd0
		x"57406d00", -- ccd4
		x"002cb07c", -- ccd8
		x"00016e00", -- ccdc
		x"0024e340", -- cce0
		x"323b0006", -- cce4
		x"4efb1002", -- cce8
		x"0004000e", -- ccec
		x"3d6effd0", -- ccf0
		x"fff06000", -- ccf4
		x"00123d6e", -- ccf8
		x"ffd2fff0", -- ccfc
		x"60000008", -- cd00
		x"3d6effd4", -- cd04
		x"fff0206e", -- cd08
		x"ffcc217c", -- cd0c
		x"003d0900", -- cd10
		x"033a4868", -- cd14
		x"033a4eba", -- cd18
		x"85026000", -- cd1c
		x"00083d6e", -- cd20
		x"ffd4fff0", -- cd24
		x"600006fc", -- cd28
		x"558f2f2e", -- cd2c
		x"fffc206e", -- cd30
		x"ffcc4868", -- cd34
		x"033a3f3c", -- cd38
		x"00812f3c", -- cd3c
		x"00000063", -- cd40
		x"486efff4", -- cd44
		x"4ebae9a2", -- cd48
		x"301f5540", -- cd4c
		x"6d00002c", -- cd50
		x"b07c0001", -- cd54
		x"6e000024", -- cd58
		x"e340323b", -- cd5c
		x"00064efb", -- cd60
		x"1002000e", -- cd64
		x"00043d6e", -- cd68
		x"ffd0fff0", -- cd6c
		x"60000012", -- cd70
		x"3d6effd2", -- cd74
		x"fff06000", -- cd78
		x"00083d6e", -- cd7c
		x"ffd4fff0", -- cd80
		x"600006a0", -- cd84
		x"2d6efff4", -- cd88
		x"ffc4206e", -- cd8c
		x"ffc44aa8", -- cd90
		x"000257c0", -- cd94
		x"4a280001", -- cd98
		x"57c1c200", -- cd9c
		x"6700000c", -- cda0
		x"3d6effd0", -- cda4
		x"fff06000", -- cda8
		x"0030206e", -- cdac
		x"ffc44aa8", -- cdb0
		x"00025ec0", -- cdb4
		x"4a680006", -- cdb8
		x"57c1c200", -- cdbc
		x"6700000c", -- cdc0
		x"3d6effd2", -- cdc4
		x"fff06000", -- cdc8
		x"00103d6e", -- cdcc
		x"ffd4fff0", -- cdd0
		x"2f2efffc", -- cdd4
		x"4ebae582", -- cdd8
		x"60000648", -- cddc
		x"558f2f0e", -- cde0
		x"4ebafbba", -- cde4
		x"4a1f6700", -- cde8
		x"0134526e", -- cdec
		x"ffea206e", -- cdf0
		x"ffec302e", -- cdf4
		x"ffeac1fc", -- cdf8
		x"001841f0", -- cdfc
		x"08e82d48", -- ce00
		x"ffc42d6e", -- ce04
		x"fff4ffc0", -- ce08
		x"206effc8", -- ce0c
		x"700a9068", -- ce10
		x"001e4440", -- ce14
		x"48c02d40", -- ce18
		x"ffde4aae", -- ce1c
		x"ffde6f00", -- ce20
		x"0010226e", -- ce24
		x"ffc07000", -- ce28
		x"1029000a", -- ce2c
		x"2d40ffde", -- ce30
		x"206effc8", -- ce34
		x"226effc4", -- ce38
		x"4ca81c00", -- ce3c
		x"000e4891", -- ce40
		x"1c004269", -- ce44
		x"0014246e", -- ce48
		x"ffc04a6a", -- ce4c
		x"00066600", -- ce50
		x"00644aae", -- ce54
		x"ffde6600", -- ce58
		x"001847fa", -- ce5c
		x"062a101b", -- ce60
		x"49e90006", -- ce64
		x"18c018db", -- ce68
		x"530062fa", -- ce6c
		x"60000016", -- ce70
		x"700db0ae", -- ce74
		x"ffde6c00", -- ce78
		x"000c206e", -- ce7c
		x"ffc0117c", -- ce80
		x"ff0d000a", -- ce84
		x"206effc0", -- ce88
		x"43e8000a", -- ce8c
		x"1019266e", -- ce90
		x"ffc445eb", -- ce94
		x"000614c0", -- ce98
		x"14d95300", -- ce9c
		x"62fa422b", -- cea0
		x"00163d6e", -- cea4
		x"ffd4fff0", -- cea8
		x"2f2efffc", -- ceac
		x"4ebae4aa", -- ceb0
		x"60000066", -- ceb4
		x"206effc4", -- ceb8
		x"117cff01", -- cebc
		x"00164aae", -- cec0
		x"ffde6f00", -- cec4
		x"00461d7c", -- cec8
		x"0001ffd9", -- cecc
		x"43fa05b8", -- ced0
		x"101945e8", -- ced4
		x"000614c0", -- ced8
		x"14d95300", -- cedc
		x"62fa226e", -- cee0
		x"ffc0246e", -- cee4
		x"ffc83569", -- cee8
		x"00060014", -- ceec
		x"3d6effd2", -- cef0
		x"fff0266e", -- cef4
		x"ffcc7000", -- cef8
		x"102b005f", -- cefc
		x"3d40ffe8", -- cf00
		x"176effeb", -- cf04
		x"005f6000", -- cf08
		x"00103d6e", -- cf0c
		x"ffd0fff0", -- cf10
		x"2f2efffc", -- cf14
		x"4ebae442", -- cf18
		x"60000010", -- cf1c
		x"3d6effd0", -- cf20
		x"fff02f2e", -- cf24
		x"fffc4eba", -- cf28
		x"e4306000", -- cf2c
		x"04f62d7c", -- cf30
		x"00002710", -- cf34
		x"ffe4486e", -- cf38
		x"ffe44eba", -- cf3c
		x"82de558f", -- cf40
		x"2f2efffc", -- cf44
		x"486effe4", -- cf48
		x"3f3c0081", -- cf4c
		x"2f3c0000", -- cf50
		x"0063486e", -- cf54
		x"fff44eba", -- cf58
		x"e790301f", -- cf5c
		x"e340323b", -- cf60
		x"00064efb", -- cf64
		x"1002001c", -- cf68
		x"00380012", -- cf6c
		x"00083d6e", -- cf70
		x"ffd0fff0", -- cf74
		x"60000028", -- cf78
		x"3d6effd2", -- cf7c
		x"fff06000", -- cf80
		x"001e4a6e", -- cf84
		x"ffe26f00", -- cf88
		x"000c3d6e", -- cf8c
		x"ffd4fff0", -- cf90
		x"60000008", -- cf94
		x"3d6effd2", -- cf98
		x"fff06000", -- cf9c
		x"00026000", -- cfa0
		x"0482206e", -- cfa4
		x"ffcc7000", -- cfa8
		x"1028005f", -- cfac
		x"b06effea", -- cfb0
		x"6d00000c", -- cfb4
		x"3d6effd2", -- cfb8
		x"fff06000", -- cfbc
		x"0034206e", -- cfc0
		x"ffcc7000", -- cfc4
		x"1028005f", -- cfc8
		x"52401140", -- cfcc
		x"005f3d7c", -- cfd0
		x"0003fff2", -- cfd4
		x"226effec", -- cfd8
		x"70001028", -- cfdc
		x"005fc1fc", -- cfe0
		x"00184a31", -- cfe4
		x"08fe6600", -- cfe8
		x"00083d6e", -- cfec
		x"ffd0fff0", -- cff0
		x"60000430", -- cff4
		x"558f486e", -- cff8
		x"fff24eba", -- cffc
		x"07664a1f", -- d000
		x"670000b6", -- d004
		x"206effec", -- d008
		x"226effcc", -- d00c
		x"70001029", -- d010
		x"005fc1fc", -- d014
		x"001841f0", -- d018
		x"08e82d48", -- d01c
		x"ffc4206e", -- d020
		x"ffc44c90", -- d024
		x"1c004891", -- d028
		x"1c0045e8", -- d02c
		x"0006101a", -- d030
		x"47e900ce", -- d034
		x"16c016da", -- d038
		x"530062fa", -- d03c
		x"30280014", -- d040
		x"5240246e", -- d044
		x"ffc848c0", -- d048
		x"25400016", -- d04c
		x"357cffff", -- d050
		x"0014558f", -- d054
		x"2f0e4eba", -- d058
		x"f9c4301f", -- d05c
		x"57406d00", -- d060
		x"003eb07c", -- d064
		x"00016e00", -- d068
		x"0036e340", -- d06c
		x"323b0006", -- d070
		x"4efb1002", -- d074
		x"0004000e", -- d078
		x"3d6effd0", -- d07c
		x"fff06000", -- d080
		x"00244a6e", -- d084
		x"ffe26f00", -- d088
		x"000c3d6e", -- d08c
		x"ffd2fff0", -- d090
		x"60000008", -- d094
		x"3d6effd0", -- d098
		x"fff06000", -- d09c
		x"00083d6e", -- d0a0
		x"ffd4fff0", -- d0a4
		x"2d7c003d", -- d0a8
		x"0900ffe4", -- d0ac
		x"486effe4", -- d0b0
		x"4eba8168", -- d0b4
		x"60000008", -- d0b8
		x"3d6effd4", -- d0bc
		x"fff06000", -- d0c0
		x"0362558f", -- d0c4
		x"2f2efffc", -- d0c8
		x"486effe4", -- d0cc
		x"3f3c0081", -- d0d0
		x"2f3c0000", -- d0d4
		x"0063486e", -- d0d8
		x"fff44eba", -- d0dc
		x"e60c301f", -- d0e0
		x"e340323b", -- d0e4
		x"00064efb", -- d0e8
		x"1002001c", -- d0ec
		x"00380012", -- d0f0
		x"00083d6e", -- d0f4
		x"ffd0fff0", -- d0f8
		x"60000028", -- d0fc
		x"3d6effd2", -- d100
		x"fff06000", -- d104
		x"001e4a6e", -- d108
		x"ffe26f00", -- d10c
		x"000c3d6e", -- d110
		x"ffd4fff0", -- d114
		x"60000008", -- d118
		x"3d6effd2", -- d11c
		x"fff06000", -- d120
		x"00026000", -- d124
		x"02fe2d6e", -- d128
		x"fff4ffc4", -- d12c
		x"206effec", -- d130
		x"226effcc", -- d134
		x"70001029", -- d138
		x"005fc1fc", -- d13c
		x"001841f0", -- d140
		x"08e82d48", -- d144
		x"ffc0206e", -- d148
		x"ffc03028", -- d14c
		x"00145240", -- d150
		x"246effc4", -- d154
		x"48c0b0aa", -- d158
		x"000256c0", -- d15c
		x"266effc8", -- d160
		x"49eb000e", -- d164
		x"7406b10c", -- d168
		x"6600000a", -- d16c
		x"538266f6", -- d170
		x"60000006", -- d174
		x"72016002", -- d178
		x"42818001", -- d17c
		x"67000014", -- d180
		x"3d6effd4", -- d184
		x"fff02f2e", -- d188
		x"fffc4eba", -- d18c
		x"e1cc6000", -- d190
		x"0028206e", -- d194
		x"ffc8317c", -- d198
		x"00070026", -- d19c
		x"226effc4", -- d1a0
		x"4a290001", -- d1a4
		x"6600000c", -- d1a8
		x"3d6effd0", -- d1ac
		x"fff06000", -- d1b0
		x"00083d6e", -- d1b4
		x"ffd2fff0", -- d1b8
		x"60000268", -- d1bc
		x"2d6efff4", -- d1c0
		x"ffc4206e", -- d1c4
		x"ffc8700a", -- d1c8
		x"9068001e", -- d1cc
		x"444048c0", -- d1d0
		x"2d40ffde", -- d1d4
		x"226effc4", -- d1d8
		x"45e9000a", -- d1dc
		x"101a286e", -- d1e0
		x"000847d4", -- d1e4
		x"16c016da", -- d1e8
		x"530062fa", -- d1ec
		x"246effcc", -- d1f0
		x"26680022", -- d1f4
		x"26aa005e", -- d1f8
		x"26680022", -- d1fc
		x"177c0000", -- d200
		x"0003266e", -- d204
		x"ffec7000", -- d208
		x"102a005f", -- d20c
		x"c1fc0018", -- d210
		x"47f308e8", -- d214
		x"2d4bffc0", -- d218
		x"266effc0", -- d21c
		x"37690004", -- d220
		x"001449eb", -- d224
		x"0006101c", -- d228
		x"47ea00ce", -- d22c
		x"16c016dc", -- d230
		x"530062fa", -- d234
		x"2f2efffc", -- d238
		x"4ebae11e", -- d23c
		x"206effc8", -- d240
		x"226effcc", -- d244
		x"4ca81c00", -- d248
		x"000e4891", -- d24c
		x"1c004229", -- d250
		x"033e4a2e", -- d254
		x"ffd96700", -- d258
		x"005a558f", -- d25c
		x"2f2efffc", -- d260
		x"4ebaf314", -- d264
		x"301f48c0", -- d268
		x"2d40ffda", -- d26c
		x"7004b0ae", -- d270
		x"ffda57c0", -- d274
		x"4aaeffda", -- d278
		x"57c18200", -- d27c
		x"67000014", -- d280
		x"4a6effe2", -- d284
		x"5ec0206e", -- d288
		x"ffcc0200", -- d28c
		x"ff011140", -- d290
		x"033e206e", -- d294
		x"ffcc4a28", -- d298
		x"033e6700", -- d29c
		x"000c226e", -- d2a0
		x"ffc8336e", -- d2a4
		x"ffd60026", -- d2a8
		x"206effcc", -- d2ac
		x"116effe9", -- d2b0
		x"005f426e", -- d2b4
		x"fff06000", -- d2b8
		x"016a2d6e", -- d2bc
		x"fff4ffc4", -- d2c0
		x"206effc4", -- d2c4
		x"7012b028", -- d2c8
		x"00016600", -- d2cc
		x"0024226e", -- d2d0
		x"ffec246e", -- d2d4
		x"ffcc7000", -- d2d8
		x"102a005f", -- d2dc
		x"c1fc0018", -- d2e0
		x"13bc0001", -- d2e4
		x"08fe3d6e", -- d2e8
		x"ffd0fff0", -- d2ec
		x"60000038", -- d2f0
		x"206effc4", -- d2f4
		x"7004b028", -- d2f8
		x"00016600", -- d2fc
		x"000c3d6e", -- d300
		x"ffd0fff0", -- d304
		x"60000020", -- d308
		x"206effc4", -- d30c
		x"7003b028", -- d310
		x"00016600", -- d314
		x"000c3d6e", -- d318
		x"ffd2fff0", -- d31c
		x"60000008", -- d320
		x"3d6effd4", -- d324
		x"fff02f2e", -- d328
		x"fffc4eba", -- d32c
		x"e02c6000", -- d330
		x"00f2206e", -- d334
		x"ffcc226e", -- d338
		x"ffc82469", -- d33c
		x"002224a8", -- d340
		x"005e2469", -- d344
		x"0022157c", -- d348
		x"00000003", -- d34c
		x"246effec", -- d350
		x"70001028", -- d354
		x"005fc1fc", -- d358
		x"001845f2", -- d35c
		x"08e82d4a", -- d360
		x"ffc4246e", -- d364
		x"ffc447ea", -- d368
		x"0006101b", -- d36c
		x"49e800ce", -- d370
		x"18c018db", -- d374
		x"530062fa", -- d378
		x"157c0001", -- d37c
		x"001645fa", -- d380
		x"010e101a", -- d384
		x"286e0008", -- d388
		x"47d416c0", -- d38c
		x"16da5300", -- d390
		x"62fa336e", -- d394
		x"ffd00026", -- d398
		x"117cff00", -- d39c
		x"005f426e", -- d3a0
		x"fff06000", -- d3a4
		x"007e422e", -- d3a8
		x"000c206e", -- d3ac
		x"ffc8316e", -- d3b0
		x"ffd00026", -- d3b4
		x"226effcc", -- d3b8
		x"137cff00", -- d3bc
		x"005f426e", -- d3c0
		x"fff06000", -- d3c4
		x"005e3d6e", -- d3c8
		x"ffd0fff0", -- d3cc
		x"2f3c000f", -- d3d0
		x"4240302e", -- d3d4
		x"ffd248c0", -- d3d8
		x"2f004eba", -- d3dc
		x"add02d5f", -- d3e0
		x"ffe4486e", -- d3e4
		x"ffe44eba", -- d3e8
		x"03566000", -- d3ec
		x"00363d6e", -- d3f0
		x"ffd0fff0", -- d3f4
		x"206effc8", -- d3f8
		x"316effd2", -- d3fc
		x"00263d6e", -- d400
		x"ffd4ffd6", -- d404
		x"6000001c", -- d408
		x"3d6effd0", -- d40c
		x"fff02f2e", -- d410
		x"fffc4eba", -- d414
		x"df446000", -- d418
		x"000a422e", -- d41c
		x"000c426e", -- d420
		x"fff04a6e", -- d424
		x"fff06600", -- d428
		x"f7ba206e", -- d42c
		x"ffc82268", -- d430
		x"001a336e", -- d434
		x"ffea0002", -- d438
		x"226effcc", -- d43c
		x"136effe3", -- d440
		x"00612b6f", -- d444
		x"0008fff6", -- d448
		x"defc000c", -- d44c
		x"4efa0032", -- d450
		x"2c5f2b5f", -- d454
		x"fff6206e", -- d458
		x"ffc82268", -- d45c
		x"001a336e", -- d460
		x"ffea0002", -- d464
		x"422e000c", -- d468
		x"7005b06d", -- d46c
		x"fffe56c0", -- d470
		x"7206b26d", -- d474
		x"fffe56c1", -- d478
		x"c2006700", -- d47c
		x"00044e4a", -- d480
		x"4e5e2e9f", -- d484
		x"4e750000", -- d488
		x"09000900", -- d48c
		x"00040f00", -- d490
		x"53657276", -- d494
		x"65722041", -- d498
		x"626f7274", -- d49c
		x"65644e75", -- d4a0
		x"60000c04", -- d4a4
		x"60000caa", -- d4a8
		x"60000cda", -- d4ac
		x"600000d6", -- d4b0
		x"4e754e75", -- d4b4
		x"2078fed4", -- d4b8
		x"43fa00da", -- d4bc
		x"21490024", -- d4c0
		x"43fa004a", -- d4c4
		x"21490028", -- d4c8
		x"4e754a90", -- d4cc
		x"670ab028", -- d4d0
		x"00086704", -- d4d4
		x"d1d060f2", -- d4d8
		x"22680004", -- d4dc
		x"4e752078", -- d4e0
		x"fed41028", -- d4e4
		x"005ec03c", -- d4e8
		x"00e02068", -- d4ec
		x"002860da", -- d4f0
		x"2078fed4", -- d4f4
		x"1028005e", -- d4f8
		x"c03c001f", -- d4fc
		x"20680024", -- d500
		x"60c861da", -- d504
		x"4ed161d6", -- d508
		x"4ee90004", -- d50c
		x"0000000a", -- d510
		x"0000d538", -- d514
		x"00000000", -- d518
		x"000a0000", -- d51c
		x"d5402000", -- d520
		x"0000000a", -- d524
		x"0000d548", -- d528
		x"40000000", -- d52c
		x"00000000", -- d530
		x"d5500000", -- d534
		x"600007c0", -- d538
		x"60000822", -- d53c
		x"60000962", -- d540
		x"600009ce", -- d544
		x"60000a70", -- d548
		x"60000ab8", -- d54c
		x"60000006", -- d550
		x"60000008", -- d554
		x"205f51d7", -- d558
		x"4ed0205f", -- d55c
		x"defc0014", -- d560
		x"51d74ed0", -- d564
		x"618a4ed1", -- d568
		x"61864ee9", -- d56c
		x"00046180", -- d570
		x"4ee90008", -- d574
		x"6100ff7a", -- d578
		x"4ee9000c", -- d57c
		x"6100ff72", -- d580
		x"4ee90010", -- d584
		x"6100ff6a", -- d588
		x"41e80009", -- d58c
		x"2f480008", -- d590
		x"4ee90004", -- d594
		x"0000000a", -- d598
		x"0000d660", -- d59c
		x"0e0f0000", -- d5a0
		x"000a0000", -- d5a4
		x"d6740f0f", -- d5a8
		x"0000000a", -- d5ac
		x"0000d638", -- d5b0
		x"040f0000", -- d5b4
		x"000a0000", -- d5b8
		x"d638050f", -- d5bc
		x"0000000a", -- d5c0
		x"0000d638", -- d5c4
		x"070f0000", -- d5c8
		x"000a0000", -- d5cc
		x"d638080f", -- d5d0
		x"0000000a", -- d5d4
		x"0000d638", -- d5d8
		x"090f0000", -- d5dc
		x"000a0000", -- d5e0
		x"d6380a2f", -- d5e4
		x"0000000a", -- d5e8
		x"0000d638", -- d5ec
		x"0b2f0000", -- d5f0
		x"000a0000", -- d5f4
		x"d6380c0f", -- d5f8
		x"0000000a", -- d5fc
		x"0000d638", -- d600
		x"0d0f0000", -- d604
		x"000a0000", -- d608
		x"d64c102f", -- d60c
		x"0000000a", -- d610
		x"0000d64c", -- d614
		x"112f0000", -- d618
		x"000a0000", -- d61c
		x"d6881609", -- d620
		x"0000000a", -- d624
		x"0000d69c", -- d628
		x"14040000", -- d62c
		x"00000000", -- d630
		x"d6b00000", -- d634
		x"60000f90", -- d638
		x"6000102a", -- d63c
		x"6000108a", -- d640
		x"600010d8", -- d644
		x"60001454", -- d648
		x"60001ae4", -- d64c
		x"60001b30", -- d650
		x"60001d0e", -- d654
		x"60001d38", -- d658
		x"60001e26", -- d65c
		x"60003a3a", -- d660
		x"6000346a", -- d664
		x"60003af4", -- d668
		x"60003864", -- d66c
		x"60003330", -- d670
		x"600039d2", -- d674
		x"60003456", -- d678
		x"60003ae0", -- d67c
		x"60003684", -- d680
		x"6000331c", -- d684
		x"6000003a", -- d688
		x"60001f7a", -- d68c
		x"6000003a", -- d690
		x"60001f90", -- d694
		x"60002020", -- d698
		x"60000026", -- d69c
		x"600000a6", -- d6a0
		x"60000026", -- d6a4
		x"600028bc", -- d6a8
		x"600028be", -- d6ac
		x"60000012", -- d6b0
		x"60000016", -- d6b4
		x"60000012", -- d6b8
		x"6000000e", -- d6bc
		x"6000000a", -- d6c0
		x"205f588f", -- d6c4
		x"51d74ed0", -- d6c8
		x"3b7c0001", -- d6cc
		x"fffe4e4a", -- d6d0
		x"558f6100", -- d6d4
		x"d340301f", -- d6d8
		x"b07c0020", -- d6dc
		x"670eb07c", -- d6e0
		x"00016708", -- d6e4
		x"b07c0008", -- d6e8
		x"66de5897", -- d6ec
		x"4e7561e0", -- d6f0
		x"60002186", -- d6f4
		x"60002582", -- d6f8
		x"61d66000", -- d6fc
		x"23866000", -- d700
		x"26b261cc", -- d704
		x"600021ca", -- d708
		x"600025b8", -- d70c
		x"61c26000", -- d710
		x"25226000", -- d714
		x"283861b8", -- d718
		x"600021dc", -- d71c
		x"600025be", -- d720
		x"61ae6000", -- d724
		x"23ac6000", -- d728
		x"26be61a4", -- d72c
		x"600023f0", -- d730
		x"600026fa", -- d734
		x"60003ad2", -- d738
		x"4ef90000", -- d73c
		x"0ae44ef9", -- d740
		x"0000521e", -- d744
		x"4ef90000", -- d748
		x"44ca4ef8", -- d74c
		x"30fe205f", -- d750
		x"301f805f", -- d754
		x"3e804ed0", -- d758
		x"205f101f", -- d75c
		x"801f1e80", -- d760
		x"4ed0205f", -- d764
		x"225f4217", -- d768
		x"4a516f06", -- d76c
		x"53511ebc", -- d770
		x"00014ed0", -- d774
		x"301b0240", -- d778
		x"000fe900", -- d77c
		x"321b0201", -- d780
		x"000f8001", -- d784
		x"4e75205f", -- d788
		x"225f245f", -- d78c
		x"264ad7fc", -- d790
		x"0000c000", -- d794
		x"61de4a00", -- d798
		x"6706d7fc", -- d79c
		x"00000040", -- d7a0
		x"61d27e00", -- d7a4
		x"1e007405", -- d7a8
		x"61cade40", -- d7ac
		x"12c051ca", -- d7b0
		x"fff87406", -- d7b4
		x"61bede40", -- d7b8
		x"51cafffa", -- d7bc
		x"61b60247", -- d7c0
		x"00ffbe00", -- d7c4
		x"57d74ed0", -- d7c8
		x"4e55ff94", -- d7cc
		x"48e7fff8", -- d7d0
		x"41fa0036", -- d7d4
		x"43edff94", -- d7d8
		x"45fa009a", -- d7dc
		x"428732d8", -- d7e0
		x"b5c866fa", -- d7e4
		x"206d000c", -- d7e8
		x"4aad0008", -- d7ec
		x"66064eba", -- d7f0
		x"00846004", -- d7f4
		x"4eba0290", -- d7f8
		x"2b470010", -- d7fc
		x"4cdf1fff", -- d800
		x"4e5d2a5f", -- d804
		x"508f4ed5", -- d808
		x"00000000", -- d80c
		x"00000000", -- d810
		x"00000000", -- d814
		x"00008018", -- d818
		x"00008020", -- d81c
		x"00008048", -- d820
		x"8000ffe0", -- d824
		x"00008028", -- d828
		x"83000000", -- d82c
		x"00000000", -- d830
		x"00000000", -- d834
		x"00010203", -- d838
		x"04050607", -- d83c
		x"08090a0b", -- d840
		x"0c0d0e0f", -- d844
		x"11121314", -- d848
		x"15160000", -- d84c
		x"00000000", -- d850
		x"00000000", -- d854
		x"00000000", -- d858
		x"00000000", -- d85c
		x"00000000", -- d860
		x"00000000", -- d864
		x"00000000", -- d868
		x"00000000", -- d86c
		x"00000000", -- d870
		x"00000000", -- d874
		x"6100003a", -- d878
		x"48e700b4", -- d87c
		x"2a7c0000", -- d880
		x"8000dbc8", -- d884
		x"43ed4000", -- d888
		x"4eb90000", -- d88c
		x"4f8e4cdf", -- d890
		x"2d002e3c", -- d894
		x"0000000e", -- d898
		x"4a00660c", -- d89c
		x"117c0001", -- d8a0
		x"00016100", -- d8a4
		x"01164287", -- d8a8
		x"117c0001", -- d8ac
		x"00014e75", -- d8b0
		x"4dfa0102", -- d8b4
		x"22482448", -- d8b8
		x"2648d3fc", -- d8bc
		x"0000c000", -- d8c0
		x"d4fc4002", -- d8c4
		x"d6fc4000", -- d8c8
		x"7e01117c", -- d8cc
		x"00000003", -- d8d0
		x"18280003", -- d8d4
		x"02040088", -- d8d8
		x"660000da", -- d8dc
		x"5287117c", -- d8e0
		x"00080003", -- d8e4
		x"18280003", -- d8e8
		x"02040008", -- d8ec
		x"670000c6", -- d8f0
		x"52876100", -- d8f4
		x"023c0804", -- d8f8
		x"00006600", -- d8fc
		x"00b85287", -- d900
		x"18280003", -- d904
		x"0204000c", -- d908
		x"0c04000c", -- d90c
		x"660000a6", -- d910
		x"52873813", -- d914
		x"0c440004", -- d918
		x"6600009a", -- d91c
		x"36bc0002", -- d920
		x"52872807", -- d924
		x"30bc0001", -- d928
		x"52875287", -- d92c
		x"18280003", -- d930
		x"020400cc", -- d934
		x"6600007e", -- d938
		x"52870c53", -- d93c
		x"00046600", -- d940
		x"00747c03", -- d944
		x"52873486", -- d948
		x"bc526600", -- d94c
		x"006851ce", -- d950
		x"fff65287", -- d954
		x"34bc0001", -- d958
		x"36bc0000", -- d95c
		x"0c530000", -- d960
		x"66000052", -- d964
		x"36bcfffe", -- d968
		x"0c53fffe", -- d96c
		x"66465287", -- d970
		x"34bc0002", -- d974
		x"36bc00ff", -- d978
		x"3c130246", -- d97c
		x"00ff0c46", -- d980
		x"00ff6630", -- d984
		x"36bc0000", -- d988
		x"3c130246", -- d98c
		x"00ff6624", -- d990
		x"528734bc", -- d994
		x"000336bc", -- d998
		x"00073c13", -- d99c
		x"02460007", -- d9a0
		x"0c460007", -- d9a4
		x"660e36bc", -- d9a8
		x"00003c13", -- d9ac
		x"02460007", -- d9b0
		x"66024e75", -- d9b4
		x"588f6000", -- d9b8
		x"fef03b7c", -- d9bc
		x"000ffffa", -- d9c0
		x"7e122b7c", -- d9c4
		x"02142536", -- d9c8
		x"ff943b7c", -- d9cc
		x"4758ff98", -- d9d0
		x"2b7c1402", -- d9d4
		x"3625ffba", -- d9d8
		x"3b7c5847", -- d9dc
		x"ffbe2b7c", -- d9e0
		x"447b9fb0", -- d9e4
		x"ffd670e4", -- d9e8
		x"72446100", -- d9ec
		x"01a00c40", -- d9f0
		x"00006600", -- d9f4
		x"008c70e0", -- d9f8
		x"724c6100", -- d9fc
		x"01900c40", -- da00
		x"00006600", -- da04
		x"007c3b7c", -- da08
		x"000dfffa", -- da0c
		x"70e4223c", -- da10
		x"00008044", -- da14
		x"3b7c5104", -- da18
		x"ffba6100", -- da1c
		x"01700c40", -- da20
		x"0000665c", -- da24
		x"70e0724c", -- da28
		x"08ed0003", -- da2c
		x"ff9b2b7c", -- da30
		x"aa68db66", -- da34
		x"ffd66100", -- da38
		x"01540c40", -- da3c
		x"00006640", -- da40
		x"70e47244", -- da44
		x"08ad0003", -- da48
		x"ff9b2b7c", -- da4c
		x"ffffffff", -- da50
		x"ffba3b7c", -- da54
		x"ffffffbe", -- da58
		x"61000132", -- da5c
		x"0c400000", -- da60
		x"661e70e4", -- da64
		x"7254243c", -- da68
		x"000668a0", -- da6c
		x"52876100", -- da70
		x"015a0806", -- da74
		x"000a6708", -- da78
		x"0804000f", -- da7c
		x"66024e75", -- da80
		x"588f6000", -- da84
		x"fe242248", -- da88
		x"24482648", -- da8c
		x"d3fc0000", -- da90
		x"c000d4fc", -- da94
		x"4002d6fc", -- da98
		x"40003b7c", -- da9c
		x"000dfffa", -- daa0
		x"610001f0", -- daa4
		x"76067e19", -- daa8
		x"720470e4", -- daac
		x"243c0006", -- dab0
		x"68a06100", -- dab4
		x"01165343", -- dab8
		x"67044a40", -- dabc
		x"66ea0c47", -- dac0
		x"0012675a", -- dac4
		x"0806000a", -- dac8
		x"66545287", -- dacc
		x"2204c27c", -- dad0
		x"03000c41", -- dad4
		x"01006746", -- dad8
		x"52872204", -- dadc
		x"c27c0700", -- dae0
		x"0c410300", -- dae4
		x"67385287", -- dae8
		x"2205c27c", -- daec
		x"1400662e", -- daf0
		x"52872204", -- daf4
		x"02414800", -- daf8
		x"0c410000", -- dafc
		x"66205287", -- db00
		x"0805000e", -- db04
		x"66185287", -- db08
		x"02860000", -- db0c
		x"dc00660e", -- db10
		x"52874a40", -- db14
		x"66080804", -- db18
		x"000d660a", -- db1c
		x"4287117c", -- db20
		x"00010001", -- db24
		x"4e754a43", -- db28
		x"6600ff7c", -- db2c
		x"7e2360ee", -- db30
		x"42847a0a", -- db34
		x"34bc0000", -- db38
		x"53856b00", -- db3c
		x"00160828", -- db40
		x"00020003", -- db44
		x"67ee36bc", -- db48
		x"00040c53", -- db4c
		x"00046604", -- db50
		x"4e757e22", -- db54
		x"78014e75", -- db58
		x"2849d2fc", -- db5c
		x"0028d8fc", -- db60
		x"0048b949", -- db64
		x"56c8fffc", -- db68
		x"4e7534bc", -- db6c
		x"000136bc", -- db70
		x"800034bc", -- db74
		x"000236bc", -- db78
		x"000034bc", -- db7c
		x"000336bc", -- db80
		x"000434bc", -- db84
		x"000036bc", -- db88
		x"004b4e75", -- db8c
		x"243c0000", -- db90
		x"27105287", -- db94
		x"61000034", -- db98
		x"0c400000", -- db9c
		x"66000028", -- dba0
		x"0804000f", -- dba4
		x"66000020", -- dba8
		x"0805000e", -- dbac
		x"66000018", -- dbb0
		x"2248d3fc", -- dbb4
		x"00008000", -- dbb8
		x"3c290022", -- dbbc
		x"0806000e", -- dbc0
		x"66000004", -- dbc4
		x"4e757001", -- dbc8
		x"4e756100", -- dbcc
		x"00940804", -- dbd0
		x"00006600", -- dbd4
		x"007e6192", -- dbd8
		x"2248d3fc", -- dbdc
		x"00008000", -- dbe0
		x"2b42fffc", -- dbe4
		x"486dfffc", -- dbe8
		x"4eb90000", -- dbec
		x"521e3813", -- dbf0
		x"08280002", -- dbf4
		x"0003660e", -- dbf8
		x"486dfffc", -- dbfc
		x"4eb90000", -- dc00
		x"523e6aea", -- dc04
		x"604c0804", -- dc08
		x"000867ec", -- dc0c
		x"08280006", -- dc10
		x"0003673c", -- dc14
		x"08040009", -- dc18
		x"67de3a29", -- dc1c
		x"001a3c29", -- dc20
		x"00260806", -- dc24
		x"000a6632", -- dc28
		x"701e5380", -- dc2c
		x"6b243813", -- dc30
		x"08280002", -- dc34
		x"000367f2", -- dc38
		x"0804000a", -- dc3c
		x"660260ea", -- dc40
		x"302dfffa", -- dc44
		x"6100ff12", -- dc48
		x"6610303c", -- dc4c
		x"00004e75", -- dc50
		x"7e123a29", -- dc54
		x"001a3c29", -- dc58
		x"0026303c", -- dc5c
		x"00014e75", -- dc60
		x"117c0008", -- dc64
		x"00036100", -- dc68
		x"fec8117c", -- dc6c
		x"00000003", -- dc70
		x"2848d9fc", -- dc74
		x"00008000", -- dc78
		x"43edff94", -- dc7c
		x"38c17233", -- dc80
		x"38d951c9", -- dc84
		x"fffc223c", -- dc88
		x"00008024", -- dc8c
		x"31801800", -- dc90
		x"4e754240", -- dc94
		x"72047405", -- dc98
		x"49edffba", -- dc9c
		x"2248d3fc", -- dca0
		x"0000c000", -- dca4
		x"08290000", -- dca8
		x"00036706", -- dcac
		x"d3fc0000", -- dcb0
		x"00401031", -- dcb4
		x"1001e148", -- dcb8
		x"10311003", -- dcbc
		x"e908e848", -- dcc0
		x"588118c0", -- dcc4
		x"51caffec", -- dcc8
		x"49edffba", -- dccc
		x"43edff94", -- dcd0
		x"7402301c", -- dcd4
		x"e15832c0", -- dcd8
		x"51cafff8", -- dcdc
		x"4e754e75", -- dce0
		x"00480140", -- dce4
		x"7f427f40", -- dce8
		x"7f430000", -- dcec
		x"00000000", -- dcf0
		x"00004e75", -- dcf4
		x"00004e56", -- dcf8
		x"fffc0c79", -- dcfc
		x"8000ffff", -- dd00
		x"fdd257c0", -- dd04
		x"0c791000", -- dd08
		x"fffffdde", -- dd0c
		x"57c1c200", -- dd10
		x"4a79ffff", -- dd14
		x"fde057c0", -- dd18
		x"c0014a79", -- dd1c
		x"fffffde8", -- dd20
		x"57c1c200", -- dd24
		x"6700002c", -- dd28
		x"1d7c0001", -- dd2c
		x"00082d79", -- dd30
		x"fffffed4", -- dd34
		x"fffc206e", -- dd38
		x"fffc2179", -- dd3c
		x"fffffdda", -- dd40
		x"00622179", -- dd44
		x"fffffde2", -- dd48
		x"006642a8", -- dd4c
		x"006a6000", -- dd50
		x"0006422e", -- dd54
		x"00084e5e", -- dd58
		x"4e750000", -- dd5c
		x"4e56fff6", -- dd60
		x"422effff", -- dd64
		x"2d79ffff", -- dd68
		x"fed4fffa", -- dd6c
		x"206efffa", -- dd70
		x"4aa80066", -- dd74
		x"5ec0122e", -- dd78
		x"ffff0841", -- dd7c
		x"0000c200", -- dd80
		x"6700010a", -- dd84
		x"4879ffff", -- dd88
		x"fdd22f3c", -- dd8c
		x"00000100", -- dd90
		x"2f280062", -- dd94
		x"4ebaf7e6", -- dd98
		x"206efffa", -- dd9c
		x"7007b0a8", -- dda0
		x"006a5cc0", -- dda4
		x"122effff", -- dda8
		x"08410000", -- ddac
		x"c2006700", -- ddb0
		x"00be2028", -- ddb4
		x"006aeb80", -- ddb8
		x"43f9ffff", -- ddbc
		x"fdd243f1", -- ddc0
		x"08002d49", -- ddc4
		x"fff6226e", -- ddc8
		x"fff63029", -- ddcc
		x"000a5240", -- ddd0
		x"6d000030", -- ddd4
		x"b07c0001", -- ddd8
		x"6e000028", -- dddc
		x"e340323b", -- dde0
		x"00064efb", -- dde4
		x"10020004", -- dde8
		x"0018217c", -- ddec
		x"00000007", -- ddf0
		x"006a217c", -- ddf4
		x"00000001", -- ddf8
		x"00666000", -- ddfc
		x"00666000", -- de00
		x"0062206e", -- de04
		x"001470ff", -- de08
		x"b05057c0", -- de0c
		x"206efff6", -- de10
		x"226e0014", -- de14
		x"3211b268", -- de18
		x"000a57c1", -- de1c
		x"82006700", -- de20
		x"0042558f", -- de24
		x"2f2e0018", -- de28
		x"48504eba", -- de2c
		x"cc164a1f", -- de30
		x"67000030", -- de34
		x"206efff6", -- de38
		x"226e0014", -- de3c
		x"32a8000a", -- de40
		x"226e0010", -- de44
		x"22a8000c", -- de48
		x"20280010", -- de4c
		x"e180226e", -- de50
		x"000c2280", -- de54
		x"226e0008", -- de58
		x"22a8001c", -- de5c
		x"1d7c0001", -- de60
		x"ffff206e", -- de64
		x"fffa52a8", -- de68
		x"006a6000", -- de6c
		x"ff2c206e", -- de70
		x"fffa7007", -- de74
		x"b0a8006a", -- de78
		x"6c00000e", -- de7c
		x"42a8006a", -- de80
		x"53a80066", -- de84
		x"52a80062", -- de88
		x"6000fee2", -- de8c
		x"1d6effff", -- de90
		x"001c4e5e", -- de94
		x"205fdefc", -- de98
		x"00144ed0", -- de9c
		x"4e750000", -- dea0
		x"4e56fff8", -- dea4
		x"0c790700", -- dea8
		x"fffffdd2", -- deac
		x"66000058", -- deb0
		x"1d7c0001", -- deb4
		x"00082d79", -- deb8
		x"fffffed4", -- debc
		x"fff82039", -- dec0
		x"fffffdee", -- dec4
		x"6c06d0bc", -- dec8
		x"000000ff", -- decc
		x"e0802d40", -- ded0
		x"fffc2f2e", -- ded4
		x"fffc2f39", -- ded8
		x"fffffdf2", -- dedc
		x"4ebaa2ce", -- dee0
		x"206efff8", -- dee4
		x"215f0062", -- dee8
		x"2f2efffc", -- deec
		x"2f39ffff", -- def0
		x"fdf64eba", -- def4
		x"a2b8206e", -- def8
		x"fff8215f", -- defc
		x"006642a8", -- df00
		x"006a6000", -- df04
		x"0006422e", -- df08
		x"00084e5e", -- df0c
		x"4e750000", -- df10
		x"4e56fffc", -- df14
		x"422e001c", -- df18
		x"2d79ffff", -- df1c
		x"fed4fffc", -- df20
		x"206efffc", -- df24
		x"4aa80066", -- df28
		x"5ec04aa8", -- df2c
		x"006a57c1", -- df30
		x"c2006700", -- df34
		x"0074217c", -- df38
		x"00000001", -- df3c
		x"006a4879", -- df40
		x"fffffdd2", -- df44
		x"2f3c0000", -- df48
		x"01002f28", -- df4c
		x"00624eba", -- df50
		x"f62c0c79", -- df54
		x"e942ffff", -- df58
		x"fdd26600", -- df5c
		x"004c41f9", -- df60
		x"fffffdd8", -- df64
		x"1018246e", -- df68
		x"001843d2", -- df6c
		x"12c012d8", -- df70
		x"530062fa", -- df74
		x"206e0014", -- df78
		x"30bce942", -- df7c
		x"206efffc", -- df80
		x"20280062", -- df84
		x"5280226e", -- df88
		x"00102280", -- df8c
		x"20280066", -- df90
		x"5380226e", -- df94
		x"000c2280", -- df98
		x"226e0008", -- df9c
		x"22b9ffff", -- dfa0
		x"fdd41d7c", -- dfa4
		x"ff01001c", -- dfa8
		x"4e5e205f", -- dfac
		x"defc0014", -- dfb0
		x"4ed04e75", -- dfb4
		x"00004e56", -- dfb8
		x"fffc0c79", -- dfbc
		x"3000ffff", -- dfc0
		x"fdd26600", -- dfc4
		x"00341d7c", -- dfc8
		x"00010008", -- dfcc
		x"2d79ffff", -- dfd0
		x"fed4fffc", -- dfd4
		x"206efffc", -- dfd8
		x"2179ffff", -- dfdc
		x"fdde0062", -- dfe0
		x"2179ffff", -- dfe4
		x"fde20066", -- dfe8
		x"42a8006a", -- dfec
		x"2179ffff", -- dff0
		x"fdd6006e", -- dff4
		x"60000006", -- dff8
		x"422e0008", -- dffc
		x"4e5e4e75", -- e000
		x"00004e56", -- e004
		x"fffc2d79", -- e008
		x"fffffed4", -- e00c
		x"fffc206e", -- e010
		x"fffc0ca8", -- e014
		x"ffffe942", -- e018
		x"006e57c0", -- e01c
		x"4aa80066", -- e020
		x"5ec1c200", -- e024
		x"4aa8006a", -- e028
		x"57c0c001", -- e02c
		x"67000066", -- e030
		x"217c0000", -- e034
		x"0001006a", -- e038
		x"226e0014", -- e03c
		x"32bce942", -- e040
		x"226e0010", -- e044
		x"22a80062", -- e048
		x"226e000c", -- e04c
		x"22a80066", -- e050
		x"226e0008", -- e054
		x"22a8006a", -- e058
		x"4879ffff", -- e05c
		x"fdd22f3c", -- e060
		x"00000100", -- e064
		x"42a74eba", -- e068
		x"f51441f9", -- e06c
		x"fffffde6", -- e070
		x"1018246e", -- e074
		x"001843d2", -- e078
		x"12c012d8", -- e07c
		x"530062fa", -- e080
		x"206e0008", -- e084
		x"20b9ffff", -- e088
		x"fdda1d7c", -- e08c
		x"ff01001c", -- e090
		x"60000006", -- e094
		x"422e001c", -- e098
		x"4e5e205f", -- e09c
		x"defc0014", -- e0a0
		x"4ed04e75", -- e0a4
		x"00004e56", -- e0a8
		x"fffa2079", -- e0ac
		x"fffffed4", -- e0b0
		x"41e8005e", -- e0b4
		x"2d48fffa", -- e0b8
		x"2f2dfff6", -- e0bc
		x"2f0e487a", -- e0c0
		x"00642b4f", -- e0c4
		x"fff6206e", -- e0c8
		x"fffa1010", -- e0cc
		x"02800000", -- e0d0
		x"001f3d40", -- e0d4
		x"fffe4eba", -- e0d8
		x"f49c206e", -- e0dc
		x"fffa1010", -- e0e0
		x"02800000", -- e0e4
		x"001f322e", -- e0e8
		x"fffe48c1", -- e0ec
		x"b0816700", -- e0f0
		x"000a3b7c", -- e0f4
		x"0001fffe", -- e0f8
		x"4e4a4879", -- e0fc
		x"fffffdd2", -- e100
		x"2f3c0000", -- e104
		x"010042a7", -- e108
		x"4ebaf472", -- e10c
		x"558f4eba", -- e110
		x"f3f21d5f", -- e114
		x"00082b6f", -- e118
		x"0008fff6", -- e11c
		x"defc000c", -- e120
		x"4efa0024", -- e124
		x"2c5f2b5f", -- e128
		x"fff6302d", -- e12c
		x"fffe48c0", -- e130
		x"2f00487a", -- e134
		x"00164eba", -- e138
		x"a0784a1f", -- e13c
		x"66000004", -- e140
		x"4e4a422e", -- e144
		x"00084e5e", -- e148
		x"4e750002", -- e14c
		x"70000000", -- e150
		x"4e560000", -- e154
		x"558f2f2e", -- e158
		x"00142f2e", -- e15c
		x"00082079", -- e160
		x"fffffed4", -- e164
		x"4868006e", -- e168
		x"2f2e000c", -- e16c
		x"2f2e0010", -- e170
		x"4ebaf394", -- e174
		x"1d5f0018", -- e178
		x"4e5e205f", -- e17c
		x"defc0010", -- e180
		x"4ed00000", -- e184
		x"4e560000", -- e188
		x"4a2e0008", -- e18c
		x"66000010", -- e190
		x"2079ffff", -- e194
		x"fed42028", -- e198
		x"006ed1ae", -- e19c
		x"00122f2e", -- e1a0
		x"000a2f2e", -- e1a4
		x"000e2f2e", -- e1a8
		x"00124eba", -- e1ac
		x"f3d04e5e", -- e1b0
		x"205fdefc", -- e1b4
		x"000e4ed0", -- e1b8
		x"4e750000", -- e1bc
		x"00010000", -- e1c0
		x"00020003", -- e1c4
		x"00040005", -- e1c8
		x"00060007", -- e1cc
		x"00080000", -- e1d0
		x"4e56fffc", -- e1d4
		x"2079ffff", -- e1d8
		x"fed441e8", -- e1dc
		x"005e2d48", -- e1e0
		x"fffc206e", -- e1e4
		x"fffc1010", -- e1e8
		x"02800000", -- e1ec
		x"001f2f00", -- e1f0
		x"487a0034", -- e1f4
		x"4eba9fba", -- e1f8
		x"4a1f6600", -- e1fc
		x"000a3b7c", -- e200
		x"0001fffe", -- e204
		x"4e4a206e", -- e208
		x"fffc1010", -- e20c
		x"02800000", -- e210
		x"001fd080", -- e214
		x"43faffa4", -- e218
		x"d2fcfff8", -- e21c
		x"3d710800", -- e220
		x"00084e5e", -- e224
		x"4e750002", -- e228
		x"0dfc0000", -- e22c
		x"4e560000", -- e230
		x"558f4eba", -- e234
		x"ff9c301f", -- e238
		x"48c02f00", -- e23c
		x"487a000e", -- e240
		x"4eba9f6e", -- e244
		x"1d5f0008", -- e248
		x"4e5e4e75", -- e24c
		x"00020780", -- e250
		x"00004e56", -- e254
		x"0000558f", -- e258
		x"4ebaff76", -- e25c
		x"301f48c0", -- e260
		x"2f00487a", -- e264
		x"000e4eba", -- e268
		x"9f481d5f", -- e26c
		x"00084e5e", -- e270
		x"4e750002", -- e274
		x"0600004d", -- e278
		x"0002001e", -- e27c
		x"00210002", -- e280
		x"00100098", -- e284
		x"0004001f", -- e288
		x"01310004", -- e28c
		x"001f0131", -- e290
		x"0006001f", -- e294
		x"01900002", -- e298
		x"00300190", -- e29c
		x"00020030", -- e2a0
		x"03200005", -- e2a4
		x"00300320", -- e2a8
		x"00090040", -- e2ac
		x"00004e56", -- e2b0
		x"fffc558f", -- e2b4
		x"4ebaff1a", -- e2b8
		x"301fc1fc", -- e2bc
		x"000641fa", -- e2c0
		x"ffb6226e", -- e2c4
		x"000841f0", -- e2c8
		x"08004c90", -- e2cc
		x"1c004891", -- e2d0
		x"1c00558f", -- e2d4
		x"4ebafefa", -- e2d8
		x"4a5f6600", -- e2dc
		x"003e486e", -- e2e0
		x"fffc4eba", -- e2e4
		x"0136102e", -- e2e8
		x"fffee288", -- e2ec
		x"02800000", -- e2f0
		x"000f2f00", -- e2f4
		x"487a002a", -- e2f8
		x"4eba9eb6", -- e2fc
		x"4a1f6700", -- e300
		x"0010206e", -- e304
		x"0008317c", -- e308
		x"00020002", -- e30c
		x"6000000c", -- e310
		x"206e0008", -- e314
		x"317c0001", -- e318
		x"00024e5e", -- e31c
		x"2e9f4e75", -- e320
		x"00020600", -- e324
		x"00004e56", -- e328
		x"fffe3f3c", -- e32c
		x"0010486e", -- e330
		x"fffe3f3c", -- e334
		x"00014eba", -- e338
		x"f3e87000", -- e33c
		x"102efffe", -- e340
		x"3d400008", -- e344
		x"4e5e4e75", -- e348
		x"0f070f05", -- e34c
		x"00004e56", -- e350
		x"00003f3c", -- e354
		x"0008558f", -- e358
		x"4ebafef8", -- e35c
		x"7000101f", -- e360
		x"48c0d080", -- e364
		x"41faffe2", -- e368
		x"48700800", -- e36c
		x"3f3c0002", -- e370
		x"4ebaf3a4", -- e374
		x"4e5e4e75", -- e378
		x"00080302", -- e37c
		x"00081402", -- e380
		x"00080206", -- e384
		x"00080102", -- e388
		x"00080502", -- e38c
		x"000a0502", -- e390
		x"00004e56", -- e394
		x"fffc302e", -- e398
		x"000c48c0", -- e39c
		x"e58041fa", -- e3a0
		x"ffd841f0", -- e3a4
		x"08002d48", -- e3a8
		x"fffc206e", -- e3ac
		x"fffc226e", -- e3b0
		x"000812a8", -- e3b4
		x"00022279", -- e3b8
		x"fffffed4", -- e3bc
		x"246e0008", -- e3c0
		x"1029005f", -- e3c4
		x"02800000", -- e3c8
		x"000f1540", -- e3cc
		x"00013f10", -- e3d0
		x"2f2e0008", -- e3d4
		x"70001028", -- e3d8
		x"00033f00", -- e3dc
		x"4ebaf338", -- e3e0
		x"4e5e205f", -- e3e4
		x"5c4f4ed0", -- e3e8
		x"00004e56", -- e3ec
		x"fffe3f3c", -- e3f0
		x"0003486e", -- e3f4
		x"fffe4eba", -- e3f8
		x"ff9a4e5e", -- e3fc
		x"4e750000", -- e400
		x"4e560000", -- e404
		x"558f4eba", -- e408
		x"fe244a1f", -- e40c
		x"66000006", -- e410
		x"4ebaf2fa", -- e414
		x"4e5e4e75", -- e418
		x"00004e56", -- e41c
		x"fffe4267", -- e420
		x"486efffe", -- e424
		x"4ebaff6c", -- e428
		x"4ebaffd6", -- e42c
		x"3f3c0008", -- e430
		x"2f2e0008", -- e434
		x"3f3c0004", -- e438
		x"4ebaf2e6", -- e43c
		x"4e5e2e9f", -- e440
		x"4e750000", -- e444
		x"4e56ffec", -- e448
		x"486efffa", -- e44c
		x"4ebafe60", -- e450
		x"2f2e0008", -- e454
		x"302efffe", -- e458
		x"48c02f00", -- e45c
		x"4eba9d4a", -- e460
		x"201f1d40", -- e464
		x"fff52f2e", -- e468
		x"0008302e", -- e46c
		x"fffe48c0", -- e470
		x"2f004eba", -- e474
		x"9d302d5f", -- e478
		x"fff6558f", -- e47c
		x"4ebafdd4", -- e480
		x"4a1f6700", -- e484
		x"004e2079", -- e488
		x"fffffed4", -- e48c
		x"1028005f", -- e490
		x"e8880280", -- e494
		x"0000000f", -- e498
		x"e3802f2e", -- e49c
		x"fff6322e", -- e4a0
		x"fffa48c1", -- e4a4
		x"2f012d40", -- e4a8
		x"ffec4eba", -- e4ac
		x"9cf8202e", -- e4b0
		x"ffecd09f", -- e4b4
		x"1d40fff4", -- e4b8
		x"2f2efff6", -- e4bc
		x"302efffa", -- e4c0
		x"48c02f00", -- e4c4
		x"4eba9ce2", -- e4c8
		x"201f3d40", -- e4cc
		x"fff26000", -- e4d0
		x"002e2f2e", -- e4d4
		x"fff6302e", -- e4d8
		x"fffc48c0", -- e4dc
		x"2f004eba", -- e4e0
		x"9cc8201f", -- e4e4
		x"1d40fff4", -- e4e8
		x"2f2efff6", -- e4ec
		x"302efffc", -- e4f0
		x"48c02f00", -- e4f4
		x"4eba9cae", -- e4f8
		x"201f3d40", -- e4fc
		x"fff23f3c", -- e500
		x"0002486e", -- e504
		x"fff04eba", -- e508
		x"fe8a4e5e", -- e50c
		x"2e9f4e75", -- e510
		x"00004e56", -- e514
		x"fff03f3c", -- e518
		x"0001486e", -- e51c
		x"fffe4eba", -- e520
		x"fe724eba", -- e524
		x"fedc3f3c", -- e528
		x"0008486e", -- e52c
		x"fffa3f3c", -- e530
		x"00044eba", -- e534
		x"f1ec486e", -- e538
		x"fff44eba", -- e53c
		x"fd72558f", -- e540
		x"4ebafd10", -- e544
		x"4a1f6700", -- e548
		x"003c2079", -- e54c
		x"fffffed4", -- e550
		x"1028005f", -- e554
		x"e8880280", -- e558
		x"0000000f", -- e55c
		x"e3807200", -- e560
		x"122efffc", -- e564
		x"9280302e", -- e568
		x"fff448c0", -- e56c
		x"2f002f01", -- e570
		x"4eba9c3a", -- e574
		x"302efffa", -- e578
		x"48c0d09f", -- e57c
		x"2d40fff0", -- e580
		x"60000016", -- e584
		x"302efffa", -- e588
		x"c1eefff6", -- e58c
		x"7200122e", -- e590
		x"fffcd081", -- e594
		x"2d40fff0", -- e598
		x"302efff8", -- e59c
		x"48c02f00", -- e5a0
		x"2f2efff0", -- e5a4
		x"4eba9c06", -- e5a8
		x"7000102e", -- e5ac
		x"fffdd09f", -- e5b0
		x"2d400008", -- e5b4
		x"4e5e4e75", -- e5b8
		x"4e750081", -- e5bc
		x"01040106", -- e5c0
		x"010a010f", -- e5c4
		x"00004e56", -- e5c8
		x"fffc558f", -- e5cc
		x"4ebafc02", -- e5d0
		x"301f48c0", -- e5d4
		x"2f00487a", -- e5d8
		x"00504eba", -- e5dc
		x"9bd44a1f", -- e5e0
		x"67000028", -- e5e4
		x"558f4eba", -- e5e8
		x"fbe8301f", -- e5ec
		x"48c0d080", -- e5f0
		x"41faffc8", -- e5f4
		x"322e0008", -- e5f8
		x"b2700800", -- e5fc
		x"57c00200", -- e600
		x"08011d40", -- e604
		x"000c6000", -- e608
		x"0016302e", -- e60c
		x"000848c0", -- e610
		x"2f00487a", -- e614
		x"00104eba", -- e618
		x"9b981d5f", -- e61c
		x"000c4e5e", -- e620
		x"2e9f4e75", -- e624
		x"00023000", -- e628
		x"0002f800", -- e62c
		x"04393839", -- e630
		x"35200538", -- e634
		x"32393058", -- e638
		x"05393133", -- e63c
		x"58410539", -- e640
		x"31335842", -- e644
		x"05393133", -- e648
		x"58430437", -- e64c
		x"39303520", -- e650
		x"04373930", -- e654
		x"36200437", -- e658
		x"39323020", -- e65c
		x"04373932", -- e660
		x"35200000", -- e664
		x"4e56fef8", -- e668
		x"41eeff00", -- e66c
		x"43fa0054", -- e670
		x"101945d0", -- e674
		x"14c014d9", -- e678
		x"530062fa", -- e67c
		x"558f2d48", -- e680
		x"fefc4eba", -- e684
		x"fb4c206e", -- e688
		x"fefc301f", -- e68c
		x"c1fc0006", -- e690
		x"43faff9a", -- e694
		x"1f3cffff", -- e698
		x"48504871", -- e69c
		x"08002d48", -- e6a0
		x"fef84eba", -- e6a4
		x"9b24206e", -- e6a8
		x"fef843d0", -- e6ac
		x"1019246e", -- e6b0
		x"000841d2", -- e6b4
		x"10c010d9", -- e6b8
		x"530062fa", -- e6bc
		x"4e5e2e9f", -- e6c0
		x"4e750248", -- e6c4
		x"50000000", -- e6c8
		x"4e560000", -- e6cc
		x"4ebaf034", -- e6d0
		x"4ebaf03a", -- e6d4
		x"4e5e4e75", -- e6d8
		x"00004e56", -- e6dc
		x"0000558f", -- e6e0
		x"4ebac332", -- e6e4
		x"7008b05f", -- e6e8
		x"57c02079", -- e6ec
		x"fffffed4", -- e6f0
		x"08280005", -- e6f4
		x"000b56c1", -- e6f8
		x"4401c200", -- e6fc
		x"02010001", -- e700
		x"08410000", -- e704
		x"02010001", -- e708
		x"1d410008", -- e70c
		x"4e5e4e75", -- e710
		x"000b000c", -- e714
		x"000a000d", -- e718
		x"00004e56", -- e71c
		x"ffd62079", -- e720
		x"fffffed4", -- e724
		x"41e8005e", -- e728
		x"2d48fff6", -- e72c
		x"206efff6", -- e730
		x"10280001", -- e734
		x"02800000", -- e738
		x"000f7207", -- e73c
		x"b2805dc0", -- e740
		x"12280001", -- e744
		x"e8890281", -- e748
		x"0000000f", -- e74c
		x"7401b481", -- e750
		x"5dc18200", -- e754
		x"6700000a", -- e758
		x"3b7c0001", -- e75c
		x"fffe4e4a", -- e760
		x"4ebaef8c", -- e764
		x"558f4eba", -- e768
		x"ef903d5f", -- e76c
		x"fffe7003", -- e770
		x"b06efffe", -- e774
		x"57c0206e", -- e778
		x"fff61228", -- e77c
		x"00010281", -- e780
		x"0000000f", -- e784
		x"56c1558f", -- e788
		x"48ee0003", -- e78c
		x"ffee4eba", -- e790
		x"ff4a4cee", -- e794
		x"0003ffee", -- e798
		x"821fc200", -- e79c
		x"206efff6", -- e7a0
		x"7003b028", -- e7a4
		x"000155c0", -- e7a8
		x"558f48ee", -- e7ac
		x"0003ffe6", -- e7b0
		x"4ebafa7a", -- e7b4
		x"4cee0003", -- e7b8
		x"ffe6141f", -- e7bc
		x"02020001", -- e7c0
		x"08420000", -- e7c4
		x"c002558f", -- e7c8
		x"558f48ee", -- e7cc
		x"0003ffde", -- e7d0
		x"4ebac242", -- e7d4
		x"4cee0003", -- e7d8
		x"ffde3f2e", -- e7dc
		x"fffe48ee", -- e7e0
		x"0003ffd6", -- e7e4
		x"4ebafde0", -- e7e8
		x"4cee0003", -- e7ec
		x"ffd6141f", -- e7f0
		x"02020001", -- e7f4
		x"08420000", -- e7f8
		x"80028200", -- e7fc
		x"6700000a", -- e800
		x"3b7c0001", -- e804
		x"fffe4e4a", -- e808
		x"558f4eba", -- e80c
		x"fb1a4a5f", -- e810
		x"67000002", -- e814
		x"486efffa", -- e818
		x"4ebafc00", -- e81c
		x"558f4eba", -- e820
		x"fb064a5f", -- e824
		x"6700000a", -- e828
		x"3b7c0006", -- e82c
		x"fffe4e4a", -- e830
		x"102efffd", -- e834
		x"02800000", -- e838
		x"00037202", -- e83c
		x"b2806600", -- e840
		x"000a3b7c", -- e844
		x"0001fffe", -- e848
		x"4e4a558f", -- e84c
		x"4ebaf9de", -- e850
		x"4a1f6700", -- e854
		x"007a102e", -- e858
		x"fffce288", -- e85c
		x"02800000", -- e860
		x"000f2f00", -- e864
		x"487a006c", -- e868
		x"4eba9946", -- e86c
		x"4a1f6600", -- e870
		x"000a3b7c", -- e874
		x"0001fffe", -- e878
		x"4e4a102e", -- e87c
		x"fffce288", -- e880
		x"02800000", -- e884
		x"000fd080", -- e888
		x"206efff6", -- e88c
		x"43fafe82", -- e890
		x"0210fee0", -- e894
		x"30310800", -- e898
		x"81101028", -- e89c
		x"0001e888", -- e8a0
		x"02800000", -- e8a4
		x"000f56c0", -- e8a8
		x"558f2d40", -- e8ac
		x"fff24eba", -- e8b0
		x"f9a2202e", -- e8b4
		x"fff2121f", -- e8b8
		x"0201ff01", -- e8bc
		x"08410000", -- e8c0
		x"c0016700", -- e8c4
		x"000a3b7c", -- e8c8
		x"0001fffe", -- e8cc
		x"4e4a4e5e", -- e8d0
		x"4e750002", -- e8d4
		x"f0000001", -- e8d8
		x"4e56fff4", -- e8dc
		x"486efffc", -- e8e0
		x"4ebafb38", -- e8e4
		x"558f4eba", -- e8e8
		x"fa3e4a5f", -- e8ec
		x"6700000a", -- e8f0
		x"3b7c0006", -- e8f4
		x"fffe4e4a", -- e8f8
		x"102efffc", -- e8fc
		x"02800000", -- e900
		x"001f5780", -- e904
		x"6d000184", -- e908
		x"b0bc0000", -- e90c
		x"001c6e00", -- e910
		x"017ae380", -- e914
		x"323b0006", -- e918
		x"4efb1002", -- e91c
		x"00d6016e", -- e920
		x"016e016e", -- e924
		x"003a003a", -- e928
		x"003a016e", -- e92c
		x"016e003a", -- e930
		x"003a003a", -- e934
		x"003a00ca", -- e938
		x"00ca003a", -- e93c
		x"00e2016e", -- e940
		x"016e016e", -- e944
		x"00d6016e", -- e948
		x"016e016e", -- e94c
		x"016e016e", -- e950
		x"016e016e", -- e954
		x"00e2598f", -- e958
		x"4ebafbb8", -- e95c
		x"2d5ffff8", -- e960
		x"102efffc", -- e964
		x"02800000", -- e968
		x"001f7207", -- e96c
		x"b2806600", -- e970
		x"0022558f", -- e974
		x"4ebaf8b6", -- e978
		x"4a1f6700", -- e97c
		x"000e4eba", -- e980
		x"fa6a4eba", -- e984
		x"ed886000", -- e988
		x"000a3b7c", -- e98c
		x"0004fffe", -- e990
		x"4e4a206e", -- e994
		x"0008202e", -- e998
		x"fff8b0a8", -- e99c
		x"00086600", -- e9a0
		x"00245268", -- e9a4
		x"fffe700a", -- e9a8
		x"b068fffe", -- e9ac
		x"6e00000a", -- e9b0
		x"3b7c0004", -- e9b4
		x"fffe4e4a", -- e9b8
		x"206e0008", -- e9bc
		x"4228fffc", -- e9c0
		x"60000020", -- e9c4
		x"206e0008", -- e9c8
		x"317c0001", -- e9cc
		x"fffe202e", -- e9d0
		x"fff890a8", -- e9d4
		x"0008e180", -- e9d8
		x"2140fff8", -- e9dc
		x"117cff01", -- e9e0
		x"fffc6000", -- e9e4
		x"00ae3b7c", -- e9e8
		x"0004fffe", -- e9ec
		x"4e4a6000", -- e9f0
		x"00a23b7c", -- e9f4
		x"0001fffe", -- e9f8
		x"4e4a6000", -- e9fc
		x"0096082e", -- ea00
		x"0004ffff", -- ea04
		x"56c04400", -- ea08
		x"4a006700", -- ea0c
		x"000a3b7c", -- ea10
		x"0005fffe", -- ea14
		x"4e4a102e", -- ea18
		x"ffff0280", -- ea1c
		x"00000003", -- ea20
		x"67000022", -- ea24
		x"558f4eba", -- ea28
		x"f8044a1f", -- ea2c
		x"6700000e", -- ea30
		x"3b7c0003", -- ea34
		x"fffe4e4a", -- ea38
		x"6000000a", -- ea3c
		x"3b7c0002", -- ea40
		x"fffe4e4a", -- ea44
		x"206e0008", -- ea48
		x"2028000c", -- ea4c
		x"53806c06", -- ea50
		x"d0bc0000", -- ea54
		x"00ffe080", -- ea58
		x"d0a80008", -- ea5c
		x"598f2d40", -- ea60
		x"fff44eba", -- ea64
		x"faae202e", -- ea68
		x"fff4b09f", -- ea6c
		x"6c000010", -- ea70
		x"206e0008", -- ea74
		x"117c0001", -- ea78
		x"fffc6000", -- ea7c
		x"000a3b7c", -- ea80
		x"0004fffe", -- ea84
		x"4e4a6000", -- ea88
		x"000a3b7c", -- ea8c
		x"0006fffe", -- ea90
		x"4e4a4e5e", -- ea94
		x"2e9f4e75", -- ea98
		x"00004e56", -- ea9c
		x"ffe8558f", -- eaa0
		x"4ebaf78a", -- eaa4
		x"4a1f6700", -- eaa8
		x"00184eba", -- eaac
		x"f8a24eba", -- eab0
		x"ec5c558f", -- eab4
		x"4ebafc24", -- eab8
		x"1d5ffffd", -- eabc
		x"60000036", -- eac0
		x"558f4eba", -- eac4
		x"f70c7001", -- eac8
		x"b05f6600", -- eacc
		x"0024486e", -- ead0
		x"ffe84eba", -- ead4
		x"f946082e", -- ead8
		x"0000ffea", -- eadc
		x"56c04400", -- eae0
		x"08400000", -- eae4
		x"02000001", -- eae8
		x"1d40fffd", -- eaec
		x"60000006", -- eaf0
		x"422efffd", -- eaf4
		x"4a2efffd", -- eaf8
		x"67000018", -- eafc
		x"2f2e0008", -- eb00
		x"4ebaf942", -- eb04
		x"4ebaec06", -- eb08
		x"3d7c0005", -- eb0c
		x"fff26000", -- eb10
		x"00083d7c", -- eb14
		x"0004fff2", -- eb18
		x"426efffe", -- eb1c
		x"4aae000c", -- eb20
		x"6f000136", -- eb24
		x"4a2efffd", -- eb28
		x"6700000e", -- eb2c
		x"2d7c0000", -- eb30
		x"0100fff4", -- eb34
		x"6000006a", -- eb38
		x"2f2e0008", -- eb3c
		x"4ebaf906", -- eb40
		x"558f4eba", -- eb44
		x"f6e84a1f", -- eb48
		x"6700004a", -- eb4c
		x"2d7c0001", -- eb50
		x"0000fff4", -- eb54
		x"558f4eba", -- eb58
		x"f6fa4a1f", -- eb5c
		x"67000032", -- eb60
		x"202e0008", -- eb64
		x"e1802f00", -- eb68
		x"2f3c004b", -- eb6c
		x"00004eba", -- eb70
		x"9638203c", -- eb74
		x"004b0000", -- eb78
		x"909f2d40", -- eb7c
		x"ffec202e", -- eb80
		x"ffecb0ae", -- eb84
		x"fff46c00", -- eb88
		x"00082d6e", -- eb8c
		x"ffecfff4", -- eb90
		x"6000000a", -- eb94
		x"2d7c7fff", -- eb98
		x"fffffff4", -- eb9c
		x"4ebaeb6e", -- eba0
		x"202e000c", -- eba4
		x"b0aefff4", -- eba8
		x"6e00000c", -- ebac
		x"2d6e000c", -- ebb0
		x"fff86000", -- ebb4
		x"00082d6e", -- ebb8
		x"fff4fff8", -- ebbc
		x"3f2efff2", -- ebc0
		x"486efff0", -- ebc4
		x"4ebaf7cc", -- ebc8
		x"4ebaf836", -- ebcc
		x"2f2dfff6", -- ebd0
		x"2f0e487a", -- ebd4
		x"00242b4f", -- ebd8
		x"fff64267", -- ebdc
		x"2f2e0010", -- ebe0
		x"2f2efff8", -- ebe4
		x"42674eba", -- ebe8
		x"eb422b6f", -- ebec
		x"0008fff6", -- ebf0
		x"defc000c", -- ebf4
		x"4efa0014", -- ebf8
		x"2c5f2b5f", -- ebfc
		x"fff67006", -- ec00
		x"b06dfffe", -- ec04
		x"67000004", -- ec08
		x"4e4a4eba", -- ec0c
		x"eb00558f", -- ec10
		x"4ebaf714", -- ec14
		x"4a5f6600", -- ec18
		x"000c1d7c", -- ec1c
		x"0001fffc", -- ec20
		x"60000008", -- ec24
		x"2f0e4eba", -- ec28
		x"fcb04a2e", -- ec2c
		x"fffc6700", -- ec30
		x"0024202e", -- ec34
		x"fff86c06", -- ec38
		x"d0bc0000", -- ec3c
		x"00ffe080", -- ec40
		x"d1ae0008", -- ec44
		x"202efff8", -- ec48
		x"d1ae0010", -- ec4c
		x"202efff8", -- ec50
		x"91ae000c", -- ec54
		x"6000fec6", -- ec58
		x"4e5e205f", -- ec5c
		x"defc000c", -- ec60
		x"4ed04e75", -- ec64
		x"00004e56", -- ec68
		x"fffe3f3c", -- ec6c
		x"0010486e", -- ec70
		x"fffe3f3c", -- ec74
		x"00014eba", -- ec78
		x"eaa87000", -- ec7c
		x"102efffe", -- ec80
		x"3d400008", -- ec84
		x"4e5e4e75", -- ec88
		x"00004e56", -- ec8c
		x"fffe2079", -- ec90
		x"fffffed4", -- ec94
		x"1028005f", -- ec98
		x"02800000", -- ec9c
		x"000f7220", -- eca0
		x"d2801d41", -- eca4
		x"fffe1d7c", -- eca8
		x"ff08ffff", -- ecac
		x"3f3c0012", -- ecb0
		x"486efffe", -- ecb4
		x"3f3c0002", -- ecb8
		x"4ebaea5c", -- ecbc
		x"4ebaea4e", -- ecc0
		x"558f4eba", -- ecc4
		x"ffa23d5f", -- ecc8
		x"00084e5e", -- eccc
		x"4e750000", -- ecd0
		x"4e56fffe", -- ecd4
		x"1d6e0009", -- ecd8
		x"fffe3f3c", -- ecdc
		x"0005486e", -- ece0
		x"fffe3f3c", -- ece4
		x"00014eba", -- ece8
		x"ea2e4e5e", -- ecec
		x"205f544f", -- ecf0
		x"4ed00000", -- ecf4
		x"4e56fffe", -- ecf8
		x"7020d06e", -- ecfc
		x"000a1d40", -- ed00
		x"fffe1d6e", -- ed04
		x"0009ffff", -- ed08
		x"3f3c0005", -- ed0c
		x"486efffe", -- ed10
		x"3f3c0002", -- ed14
		x"4ebaea00", -- ed18
		x"4e5e2e9f", -- ed1c
		x"4e750000", -- ed20
		x"4e560000", -- ed24
		x"3f3c000d", -- ed28
		x"4ebaffa6", -- ed2c
		x"4ebae9de", -- ed30
		x"3f3c000e", -- ed34
		x"2f2e0008", -- ed38
		x"3f3c0014", -- ed3c
		x"4ebae9e2", -- ed40
		x"4ebae9ca", -- ed44
		x"558f4eba", -- ed48
		x"ff1e3d5f", -- ed4c
		x"000c4e5e", -- ed50
		x"2e9f4e75", -- ed54
		x"00004e56", -- ed58
		x"00002079", -- ed5c
		x"fffffed4", -- ed60
		x"1028005f", -- ed64
		x"02800000", -- ed68
		x"000f3f00", -- ed6c
		x"3f3c0035", -- ed70
		x"4ebaff82", -- ed74
		x"4ebae996", -- ed78
		x"3f3c000e", -- ed7c
		x"2f2e0008", -- ed80
		x"3f3c0025", -- ed84
		x"4ebae99a", -- ed88
		x"4ebae982", -- ed8c
		x"558f4eba", -- ed90
		x"fed63d5f", -- ed94
		x"000c4e5e", -- ed98
		x"2e9f4e75", -- ed9c
		x"00004e56", -- eda0
		x"00007020", -- eda4
		x"d06e0008", -- eda8
		x"3f004eba", -- edac
		x"ff244eba", -- edb0
		x"e95c558f", -- edb4
		x"4ebafeb0", -- edb8
		x"3d5f000a", -- edbc
		x"4e5e205f", -- edc0
		x"544f4ed0", -- edc4
		x"00004e56", -- edc8
		x"ffee206e", -- edcc
		x"00082d58", -- edd0
		x"fff82d50", -- edd4
		x"fffc1d7c", -- edd8
		x"ff34ffee", -- eddc
		x"1d7cff3e", -- ede0
		x"ffef4cae", -- ede4
		x"0f00fff8", -- ede8
		x"48ae0f00", -- edec
		x"fff03f3c", -- edf0
		x"0005486e", -- edf4
		x"ffee3f3c", -- edf8
		x"000a4eba", -- edfc
		x"e91a4eba", -- ee00
		x"e90c558f", -- ee04
		x"4ebafe60", -- ee08
		x"3d5f000c", -- ee0c
		x"4e5e2e9f", -- ee10
		x"4e750000", -- ee14
		x"4e56fff0", -- ee18
		x"2079ffff", -- ee1c
		x"fed41028", -- ee20
		x"005fe888", -- ee24
		x"02800000", -- ee28
		x"000f7240", -- ee2c
		x"d2801d41", -- ee30
		x"fff01d7c", -- ee34
		x"ff10fff1", -- ee38
		x"426efff2", -- ee3c
		x"2d6e000e", -- ee40
		x"fff41d7c", -- ee44
		x"0034fff8", -- ee48
		x"1d7c0018", -- ee4c
		x"fff92d6e", -- ee50
		x"000afffa", -- ee54
		x"1d6e0009", -- ee58
		x"fffe3f3c", -- ee5c
		x"0005486e", -- ee60
		x"fff03f3c", -- ee64
		x"000f4eba", -- ee68
		x"e8ae4e5e", -- ee6c
		x"205fdefc", -- ee70
		x"000a4ed0", -- ee74
		x"00004e56", -- ee78
		x"00003f2e", -- ee7c
		x"00083f3c", -- ee80
		x"000e4eba", -- ee84
		x"fe704eba", -- ee88
		x"e884558f", -- ee8c
		x"4ebafdd8", -- ee90
		x"3d5f000a", -- ee94
		x"4e5e205f", -- ee98
		x"544f4ed0", -- ee9c
		x"00004e56", -- eea0
		x"00002f2e", -- eea4
		x"0012302e", -- eea8
		x"000848c0", -- eeac
		x"d0ae000a", -- eeb0
		x"2f004267", -- eeb4
		x"4ebaff5e", -- eeb8
		x"4ebae852", -- eebc
		x"2f2dfff6", -- eec0
		x"2f0e487a", -- eec4
		x"00282b4f", -- eec8
		x"fff63f3c", -- eecc
		x"000e2f2e", -- eed0
		x"000e2f2e", -- eed4
		x"000a3f2e", -- eed8
		x"00084eba", -- eedc
		x"e84e2b6f", -- eee0
		x"0008fff6", -- eee4
		x"defc000c", -- eee8
		x"4efa0014", -- eeec
		x"2c5f2b5f", -- eef0
		x"fff67006", -- eef4
		x"b06dfffe", -- eef8
		x"67000004", -- eefc
		x"4e4a4eba", -- ef00
		x"e80c558f", -- ef04
		x"4ebafd60", -- ef08
		x"3d5f0016", -- ef0c
		x"4e5e205f", -- ef10
		x"defc000e", -- ef14
		x"4ed04e75", -- ef18
		x"00000000", -- ef1c
		x"00001fff", -- ef20
		x"00004e56", -- ef24
		x"fffe422e", -- ef28
		x"ffff558f", -- ef2c
		x"487affea", -- ef30
		x"4ebafe94", -- ef34
		x"4a5f6700", -- ef38
		x"000a486e", -- ef3c
		x"ffff4eba", -- ef40
		x"000e4a2e", -- ef44
		x"ffff66de", -- ef48
		x"4e5e4e75", -- ef4c
		x"00004e56", -- ef50
		x"ffe23d7c", -- ef54
		x"fffffffe", -- ef58
		x"206e0008", -- ef5c
		x"4210422e", -- ef60
		x"ffe4558f", -- ef64
		x"486effea", -- ef68
		x"4ebafdb6", -- ef6c
		x"4a5f6700", -- ef70
		x"000a3b7c", -- ef74
		x"0005fffe", -- ef78
		x"4e4a102e", -- ef7c
		x"ffea0280", -- ef80
		x"0000000f", -- ef84
		x"3d40ffe8", -- ef88
		x"422effe5", -- ef8c
		x"3d7c0040", -- ef90
		x"ffe6536e", -- ef94
		x"ffe6302e", -- ef98
		x"ffe63200", -- ef9c
		x"e841e349", -- efa0
		x"0240000f", -- efa4
		x"243610ec", -- efa8
		x"e1aa701f", -- efac
		x"e0aa4a82", -- efb0
		x"670000fa", -- efb4
		x"302effe6", -- efb8
		x"55406d00", -- efbc
		x"00eab07c", -- efc0
		x"003d6e00", -- efc4
		x"00e2e340", -- efc8
		x"323b0006", -- efcc
		x"4efb1002", -- efd0
		x"007c00d6", -- efd4
		x"00d600d6", -- efd8
		x"0086009a", -- efdc
		x"00d600d6", -- efe0
		x"00d600d6", -- efe4
		x"00d600d6", -- efe8
		x"00d600d6", -- efec
		x"00d600d6", -- eff0
		x"00d6007c", -- eff4
		x"00d600d6", -- eff8
		x"007c00d6", -- effc
		x"007c00d6", -- f000
		x"00b600b6", -- f004
		x"00b600d6", -- f008
		x"00a400b6", -- f00c
		x"00d600b6", -- f010
		x"00d60090", -- f014
		x"00d6009a", -- f018
		x"00d600d6", -- f01c
		x"009a009a", -- f020
		x"00d6009a", -- f024
		x"009a00d6", -- f028
		x"00d600d6", -- f02c
		x"00c200c2", -- f030
		x"00c200cc", -- f034
		x"00cc00cc", -- f038
		x"00cc00cc", -- f03c
		x"00cc00cc", -- f040
		x"00cc00cc", -- f044
		x"00cc00cc", -- f048
		x"00cc00cc", -- f04c
		x"3d7c0005", -- f050
		x"fffe6000", -- f054
		x"00583d7c", -- f058
		x"0001fffe", -- f05c
		x"6000004e", -- f060
		x"3d7c0003", -- f064
		x"fffe6000", -- f068
		x"00443d7c", -- f06c
		x"0004fffe", -- f070
		x"6000003a", -- f074
		x"1d7c0001", -- f078
		x"ffe4206e", -- f07c
		x"000810bc", -- f080
		x"00016000", -- f084
		x"0028206e", -- f088
		x"000810bc", -- f08c
		x"00016000", -- f090
		x"001c1d7c", -- f094
		x"0001ffe5", -- f098
		x"60000012", -- f09c
		x"1d7c0001", -- f0a0
		x"ffe46000", -- f0a4
		x"00083d7c", -- f0a8
		x"0006fffe", -- f0ac
		x"0c6e0000", -- f0b0
		x"ffe66e00", -- f0b4
		x"fede4a6e", -- f0b8
		x"fffe6d00", -- f0bc
		x"000a3b6e", -- f0c0
		x"fffefffe", -- f0c4
		x"4e4a4a2e", -- f0c8
		x"ffe56700", -- f0cc
		x"003e3d7c", -- f0d0
		x"0001ffe2", -- f0d4
		x"7006b06e", -- f0d8
		x"ffe25cc0", -- f0dc
		x"322effe2", -- f0e0
		x"4a3610f3", -- f0e4
		x"5cc1c200", -- f0e8
		x"67000020", -- f0ec
		x"558f302e", -- f0f0
		x"ffe21036", -- f0f4
		x"00f34880", -- f0f8
		x"3f004eba", -- f0fc
		x"fd7a4a5f", -- f100
		x"67000002", -- f104
		x"526effe2", -- f108
		x"60ca558f", -- f10c
		x"3f2effe8", -- f110
		x"4ebafc8c", -- f114
		x"4a5f6600", -- f118
		x"fe4a4a2e", -- f11c
		x"ffe46700", -- f120
		x"00064eba", -- f124
		x"fdfe4e5e", -- f128
		x"2e9f4e75", -- f12c
		x"00004e56", -- f130
		x"0000302e", -- f134
		x"00086c04", -- f138
		x"d07c00ff", -- f13c
		x"e0407202", -- f140
		x"b24057c0", -- f144
		x"02000001", -- f148
		x"1d40000c", -- f14c
		x"4e5e2e9f", -- f150
		x"4e750000", -- f154
		x"4e560000", -- f158
		x"558f4eba", -- f15c
		x"e59c301f", -- f160
		x"6c04d07c", -- f164
		x"00ffe040", -- f168
		x"7202b240", -- f16c
		x"6700000a", -- f170
		x"3b7c0001", -- f174
		x"fffe4e4a", -- f178
		x"4e5e4e75", -- f17c
		x"00004e56", -- f180
		x"fecc4eba", -- f184
		x"ffd0422e", -- f188
		x"ffff558f", -- f18c
		x"486effda", -- f190
		x"4ebafbc4", -- f194
		x"4a5f6700", -- f198
		x"000a486e", -- f19c
		x"ffff4eba", -- f1a0
		x"fdae4a2e", -- f1a4
		x"ffff66de", -- f1a8
		x"202effe0", -- f1ac
		x"02ae0000", -- f1b0
		x"00ffffd6", -- f1b4
		x"0280ffff", -- f1b8
		x"ff0081ae", -- f1bc
		x"ffd6422e", -- f1c0
		x"ffd141fa", -- f1c4
		x"01841018", -- f1c8
		x"246e0008", -- f1cc
		x"43d212c0", -- f1d0
		x"12d85300", -- f1d4
		x"62fa426e", -- f1d8
		x"ffd2526e", -- f1dc
		x"ffd2302e", -- f1e0
		x"ffd248c0", -- f1e4
		x"e580d0bc", -- f1e8
		x"0000000c", -- f1ec
		x"2200e881", -- f1f0
		x"e3890280", -- f1f4
		x"0000000f", -- f1f8
		x"243618d4", -- f1fc
		x"e1aa701c", -- f200
		x"e0aa3d42", -- f204
		x"ffd44a6e", -- f208
		x"ffd46700", -- f20c
		x"00081d7c", -- f210
		x"0001ffd1", -- f214
		x"4a2effd1", -- f218
		x"67000028", -- f21c
		x"206e0008", -- f220
		x"70001010", -- f224
		x"5240206e", -- f228
		x"00081080", -- f22c
		x"7030d06e", -- f230
		x"ffd4206e", -- f234
		x"0008226e", -- f238
		x"00087200", -- f23c
		x"12111180", -- f240
		x"10000c6e", -- f244
		x"0005ffd2", -- f248
		x"6d907001", -- f24c
		x"b02effdf", -- f250
		x"660000a8", -- f254
		x"558f486e", -- f258
		x"fff14267", -- f25c
		x"2079ffff", -- f260
		x"fed41028", -- f264
		x"005fe888", -- f268
		x"02800000", -- f26c
		x"000f3f00", -- f270
		x"4ebab746", -- f274
		x"4a1f6700", -- f278
		x"004441ee", -- f27c
		x"fed0226e", -- f280
		x"000845d1", -- f284
		x"101a43d0", -- f288
		x"12c012da", -- f28c
		x"530062fa", -- f290
		x"1f3c00ff", -- f294
		x"4850487a", -- f298
		x"00b42d48", -- f29c
		x"fecc4eba", -- f2a0
		x"8f28206e", -- f2a4
		x"fecc43d0", -- f2a8
		x"1019246e", -- f2ac
		x"000841d2", -- f2b0
		x"10c010d9", -- f2b4
		x"530062fa", -- f2b8
		x"60000040", -- f2bc
		x"41eefed0", -- f2c0
		x"226e0008", -- f2c4
		x"45d1101a", -- f2c8
		x"43d012c0", -- f2cc
		x"12da5300", -- f2d0
		x"62fa1f3c", -- f2d4
		x"00ff4850", -- f2d8
		x"487a0078", -- f2dc
		x"2d48fecc", -- f2e0
		x"4eba8ee6", -- f2e4
		x"206efecc", -- f2e8
		x"43d01019", -- f2ec
		x"246e0008", -- f2f0
		x"41d210c0", -- f2f4
		x"10d95300", -- f2f8
		x"62fa7002", -- f2fc
		x"b02effdf", -- f300
		x"66000040", -- f304
		x"41eefed0", -- f308
		x"226e0008", -- f30c
		x"45d1101a", -- f310
		x"43d012c0", -- f314
		x"12da5300", -- f318
		x"62fa1f3c", -- f31c
		x"00ff4850", -- f320
		x"487a0036", -- f324
		x"2d48fecc", -- f328
		x"4eba8e9e", -- f32c
		x"206efecc", -- f330
		x"43d01019", -- f334
		x"246e0008", -- f338
		x"41d210c0", -- f33c
		x"10d95300", -- f340
		x"62fa4e5e", -- f344
		x"2e9f4e75", -- f348
		x"02485000", -- f34c
		x"05205245", -- f350
		x"4d560520", -- f354
		x"46495844", -- f358
		x"05205441", -- f35c
		x"50450000", -- f360
		x"4e56fffe", -- f364
		x"4ebae39c", -- f368
		x"4ebae3a2", -- f36c
		x"558f4eba", -- f370
		x"f8f64a5f", -- f374
		x"67000012", -- f378
		x"486effff", -- f37c
		x"4ebafbd0", -- f380
		x"3b7c0006", -- f384
		x"fffe4e4a", -- f388
		x"4e5e4e75", -- f38c
		x"00004e56", -- f390
		x"ffd42079", -- f394
		x"fffffed4", -- f398
		x"1028005f", -- f39c
		x"02800000", -- f3a0
		x"000f720e", -- f3a4
		x"b2806c00", -- f3a8
		x"000a3b7c", -- f3ac
		x"0001fffe", -- f3b0
		x"4e4a4eba", -- f3b4
		x"e33a4eba", -- f3b8
		x"fd9c422e", -- f3bc
		x"ffff558f", -- f3c0
		x"4ebaf8c8", -- f3c4
		x"4a5f6700", -- f3c8
		x"000a486e", -- f3cc
		x"ffff4eba", -- f3d0
		x"fb7e4a2e", -- f3d4
		x"ffff66e2", -- f3d8
		x"4ebafb48", -- f3dc
		x"422effff", -- f3e0
		x"558f486e", -- f3e4
		x"ffd84eba", -- f3e8
		x"f96e4a5f", -- f3ec
		x"6700000a", -- f3f0
		x"486effff", -- f3f4
		x"4ebafb58", -- f3f8
		x"4a2effff", -- f3fc
		x"66de2079", -- f400
		x"fffffed4", -- f404
		x"41e8005e", -- f408
		x"2d48ffd4", -- f40c
		x"7000102e", -- f410
		x"ffee7200", -- f414
		x"122effef", -- f418
		x"d0411d40", -- f41c
		x"fffe558f", -- f420
		x"486efffe", -- f424
		x"4267206e", -- f428
		x"ffd41028", -- f42c
		x"0001e888", -- f430
		x"02800000", -- f434
		x"000f3f00", -- f438
		x"4ebab57e", -- f43c
		x"4a1f6600", -- f440
		x"000a3b7c", -- f444
		x"0001fffe", -- f448
		x"4e4a202e", -- f44c
		x"ffe0e188", -- f450
		x"7210e2a0", -- f454
		x"0c800000", -- f458
		x"01006600", -- f45c
		x"0012206e", -- f460
		x"ffd40210", -- f464
		x"ffe07010", -- f468
		x"81106000", -- f46c
		x"000e206e", -- f470
		x"ffd40210", -- f474
		x"ffe07011", -- f478
		x"81104e5e", -- f47c
		x"4e750000", -- f480
		x"4e56ffd0", -- f484
		x"4ebafcce", -- f488
		x"422effd1", -- f48c
		x"558f2079", -- f490
		x"fffffed4", -- f494
		x"1028005f", -- f498
		x"02800000", -- f49c
		x"000f3f00", -- f4a0
		x"4ebaf8fc", -- f4a4
		x"4a5f6700", -- f4a8
		x"000a486e", -- f4ac
		x"ffd14eba", -- f4b0
		x"fa9e4a2e", -- f4b4
		x"ffd166d0", -- f4b8
		x"2079ffff", -- f4bc
		x"fed41028", -- f4c0
		x"005e0280", -- f4c4
		x"0000001f", -- f4c8
		x"7210b280", -- f4cc
		x"6600000a", -- f4d0
		x"426efffe", -- f4d4
		x"600000ca", -- f4d8
		x"422effd1", -- f4dc
		x"558f486e", -- f4e0
		x"ffd84eba", -- f4e4
		x"f8724a5f", -- f4e8
		x"6700000a", -- f4ec
		x"486effd1", -- f4f0
		x"4ebafa5c", -- f4f4
		x"4a2effd1", -- f4f8
		x"66de202e", -- f4fc
		x"ffe0e188", -- f500
		x"7210e2a0", -- f504
		x"3d40ffd4", -- f508
		x"0c6e0100", -- f50c
		x"ffd46f00", -- f510
		x"0058302e", -- f514
		x"ffd40240", -- f518
		x"00ff4a40", -- f51c
		x"6700000a", -- f520
		x"3b7c0006", -- f524
		x"fffe4e4a", -- f528
		x"302effd4", -- f52c
		x"6c04d07c", -- f530
		x"00ffe040", -- f534
		x"3d40ffd6", -- f538
		x"2f2e0008", -- f53c
		x"302effd6", -- f540
		x"48c02f00", -- f544
		x"4eba8c62", -- f548
		x"201fe180", -- f54c
		x"3d40fffe", -- f550
		x"2f2e0008", -- f554
		x"302effd6", -- f558
		x"48c02f00", -- f55c
		x"4eba8c46", -- f560
		x"2d5f0008", -- f564
		x"6000003a", -- f568
		x"203c0000", -- f56c
		x"010081ee", -- f570
		x"ffd44840", -- f574
		x"4a406700", -- f578
		x"000a3b7c", -- f57c
		x"0006fffe", -- f580
		x"4e4a426e", -- f584
		x"fffe203c", -- f588
		x"00000100", -- f58c
		x"81eeffd4", -- f590
		x"48c02f00", -- f594
		x"2f2e0008", -- f598
		x"4eba8c12", -- f59c
		x"2d5f0008", -- f5a0
		x"426effd2", -- f5a4
		x"422effd1", -- f5a8
		x"558f2f2e", -- f5ac
		x"00082f2e", -- f5b0
		x"00102f2e", -- f5b4
		x"000c3f2e", -- f5b8
		x"fffe4eba", -- f5bc
		x"f8e24a5f", -- f5c0
		x"67000028", -- f5c4
		x"486effd1", -- f5c8
		x"4ebaf984", -- f5cc
		x"4a2effd1", -- f5d0
		x"67000018", -- f5d4
		x"526effd2", -- f5d8
		x"7003b06e", -- f5dc
		x"ffd26e00", -- f5e0
		x"000a3b7c", -- f5e4
		x"0004fffe", -- f5e8
		x"4e4a4a2e", -- f5ec
		x"ffd166b4", -- f5f0
		x"4e5e205f", -- f5f4
		x"defc000c", -- f5f8
		x"4ed04e75", -- f5fc
		x"48503938", -- f600
		x"3235392e", -- f604
		x"205f225f", -- f608
		x"49e90001", -- f60c
		x"700045fa", -- f610
		x"ffec0c12", -- f614
		x"002e6706", -- f618
		x"18da5200", -- f61c
		x"60f41280", -- f620
		x"4ed0612e", -- f624
		x"42290001", -- f628
		x"487800c8", -- f62c
		x"6100b45c", -- f630
		x"14bc0019", -- f634
		x"610001c0", -- f638
		x"720be36e", -- f63c
		x"72400829", -- f640
		x"00050005", -- f644
		x"6702e54e", -- f648
		x"615214bc", -- f64c
		x"00116000", -- f650
		x"01a6558f", -- f654
		x"6100b3be", -- f658
		x"7000301f", -- f65c
		x"0c40001e", -- f660
		x"660001e8", -- f664
		x"45e9000b", -- f668
		x"47e90009", -- f66c
		x"72001229", -- f670
		x"00056b24", -- f674
		x"2e010207", -- f678
		x"00073c07", -- f67c
		x"52077011", -- f680
		x"08010005", -- f684
		x"67025400", -- f688
		x"e1af2001", -- f68c
		x"e6080200", -- f690
		x"00037240", -- f694
		x"e1694e75", -- f698
		x"588f4e75", -- f69c
		x"14bc000b", -- f6a0
		x"16bc0001", -- f6a4
		x"e4491681", -- f6a8
		x"e54916bc", -- f6ac
		x"00241686", -- f6b0
		x"e04e1686", -- f6b4
		x"4e75619a", -- f6b8
		x"205f2a1f", -- f6bc
		x"261f7807", -- f6c0
		x"08010009", -- f6c4
		x"6606e58d", -- f6c8
		x"e0ad600c", -- f6cc
		x"08050000", -- f6d0
		x"670408c4", -- f6d4
		x"0010e28d", -- f6d8
		x"303c1fff", -- f6dc
		x"08290005", -- f6e0
		x"00056602", -- f6e4
		x"e4483c05", -- f6e8
		x"cc406606", -- f6ec
		x"3c058c40", -- f6f0
		x"60043c05", -- f6f4
		x"5346285f", -- f6f8
		x"2f0861a0", -- f6fc
		x"14bc0014", -- f700
		x"2c05ccc1", -- f704
		x"dc83bc87", -- f708
		x"6e00014c", -- f70c
		x"610000e8", -- f710
		x"7e006002", -- f714
		x"52453c05", -- f718
		x"618214bc", -- f71c
		x"001d6100", -- f720
		x"00d62c01", -- f724
		x"534640c2", -- f728
		x"007c0700", -- f72c
		x"08380001", -- f730
		x"feda6612", -- f734
		x"2f3c0002", -- f738
		x"46084857", -- f73c
		x"4eb8521e", -- f740
		x"201f6000", -- f744
		x"0006303c", -- f748
		x"4c0014bc", -- f74c
		x"00120884", -- f750
		x"0010670e", -- f754
		x"0f12671e", -- f758
		x"4a135346", -- f75c
		x"0c4600ff", -- f760
		x"6ef20f12", -- f764
		x"673018d3", -- f768
		x"53836f00", -- f76c
		x"008251ce", -- f770
		x"fff246c2", -- f774
		x"609e0912", -- f778
		x"676a0838", -- f77c
		x"0001feda", -- f780
		x"660e2f00", -- f784
		x"48574eb8", -- f788
		x"523e584f", -- f78c
		x"6ac6602a", -- f790
		x"53406ec0", -- f794
		x"60240912", -- f798
		x"66060f12", -- f79c
		x"66c46044", -- f7a0
		x"08380001", -- f7a4
		x"feda660e", -- f7a8
		x"2f004857", -- f7ac
		x"4eb8523e", -- f7b0
		x"584f6aae", -- f7b4
		x"60045340", -- f7b8
		x"6ea846c2", -- f7bc
		x"60000094", -- f7c0
		x"09126606", -- f7c4
		x"0f126620", -- f7c8
		x"601a0838", -- f7cc
		x"0001feda", -- f7d0
		x"660c2f00", -- f7d4
		x"48574eb8", -- f7d8
		x"523e584f", -- f7dc
		x"6a0a5340", -- f7e0
		x"6e0660d6", -- f7e4
		x"46c26066", -- f7e8
		x"0f1267d4", -- f7ec
		x"4a1351ce", -- f7f0
		x"fff846c2", -- f7f4
		x"4e750838", -- f7f8
		x"0001feda", -- f7fc
		x"66102f3c", -- f800
		x"0016e360", -- f804
		x"48574eb8", -- f808
		x"521e201f", -- f80c
		x"6006203c", -- f810
		x"0003a000", -- f814
		x"08120007", -- f818
		x"66080812", -- f81c
		x"00066702", -- f820
		x"4e750838", -- f824
		x"0001feda", -- f828
		x"661a2f00", -- f82c
		x"48574eb8", -- f830
		x"523e588f", -- f834
		x"6ade0812", -- f838
		x"00076616", -- f83c
		x"08120006", -- f840
		x"67104e75", -- f844
		x"53806ecc", -- f848
		x"60087001", -- f84c
		x"600a7004", -- f850
		x"60067005", -- f854
		x"60027006", -- f858
		x"3b40fffe", -- f85c
		x"2e6dfff6", -- f860
		x"4e754e75", -- f864
		x"3b40fffe", -- f868
		x"4e4a45e9", -- f86c
		x"001147e9", -- f870
		x"001749e9", -- f874
		x"001f4e75", -- f878
		x"61f07001", -- f87c
		x"08290007", -- f880
		x"000567e0", -- f884
		x"70001340", -- f888
		x"000316bc", -- f88c
		x"008014bc", -- f890
		x"00081340", -- f894
		x"00131340", -- f898
		x"001b1340", -- f89c
		x"001d1340", -- f8a0
		x"001916bc", -- f8a4
		x"000e16bc", -- f8a8
		x"009316bc", -- f8ac
		x"001616bc", -- f8b0
		x"000016bc", -- f8b4
		x"001016bc", -- f8b8
		x"008f4878", -- f8bc
		x"00646100", -- f8c0
		x"b1ca16bc", -- f8c4
		x"000f16bc", -- f8c8
		x"009016bc", -- f8cc
		x"000b4e75", -- f8d0
		x"61983f3c", -- f8d4
		x"0010614e", -- f8d8
		x"611816bc", -- f8dc
		x"000818bc", -- f8e0
		x"0000610e", -- f8e4
		x"16bc000c", -- f8e8
		x"610818bc", -- f8ec
		x"00046000", -- f8f0
		x"00746000", -- f8f4
		x"00d04e56", -- f8f8
		x"00006100", -- f8fc
		x"ff6e3f2e", -- f900
		x"000e6122", -- f904
		x"206e000a", -- f908
		x"302e0008", -- f90c
		x"61e45340", -- f910
		x"6f041898", -- f914
		x"60f616bc", -- f918
		x"00081890", -- f91c
		x"61404e5e", -- f920
		x"205f508f", -- f924
		x"4ed016bc", -- f928
		x"000c61c6", -- f92c
		x"18bc00bf", -- f930
		x"613e803c", -- f934
		x"0040615e", -- f938
		x"61b81880", -- f93c
		x"16bc008a", -- f940
		x"6148803c", -- f944
		x"0020614e", -- f948
		x"61a81880", -- f94c
		x"205f7060", -- f950
		x"805f2f08", -- f954
		x"6140615e", -- f958
		x"16bc000b", -- f95c
		x"4e756164", -- f960
		x"16bc000c", -- f964
		x"615e18bc", -- f968
		x"00bf16bc", -- f96c
		x"000b6054", -- f970
		x"7015b3fc", -- f974
		x"00478000", -- f978
		x"670e701f", -- f97c
		x"c0290005", -- f980
		x"b03c001f", -- f984
		x"66027000", -- f988
		x"4e752078", -- f98c
		x"fed47000", -- f990
		x"10280061", -- f994
		x"4e751200", -- f998
		x"1401e30a", -- f99c
		x"b5011401", -- f9a0
		x"e50ab501", -- f9a4
		x"1401e90a", -- f9a8
		x"b5010201", -- f9ac
		x"0080b300", -- f9b0
		x"0a000080", -- f9b4
		x"4e75610c", -- f9b8
		x"48780055", -- f9bc
		x"6100b0cc", -- f9c0
		x"18804e75", -- f9c4
		x"76046002", -- f9c8
		x"76051212", -- f9cc
		x"07016702", -- f9d0
		x"4e750838", -- f9d4
		x"0001feda", -- f9d8
		x"66224878", -- f9dc
		x"61a84857", -- f9e0
		x"6100dd5c", -- f9e4
		x"241f8212", -- f9e8
		x"070166e4", -- f9ec
		x"2f024857", -- f9f0
		x"6100057c", -- f9f4
		x"6aee588f", -- f9f8
		x"74006004", -- f9fc
		x"343c192b", -- fa00
		x"82120701", -- fa04
		x"56cafffa", -- fa08
		x"66c67001", -- fa0c
		x"3f006100", -- fa10
		x"fe68301f", -- fa14
		x"6000fe4e", -- fa18
		x"16bc000c", -- fa1c
		x"61a618bc", -- fa20
		x"00bf6100", -- fa24
		x"ff4c803c", -- fa28
		x"00206100", -- fa2c
		x"ff6a6194", -- fa30
		x"188016bc", -- fa34
		x"0089205f", -- fa38
		x"7040805f", -- fa3c
		x"6100ff58", -- fa40
		x"61821880", -- fa44
		x"7060805f", -- fa48
		x"6100ff4c", -- fa4c
		x"6100ff68", -- fa50
		x"6100ff72", -- fa54
		x"48780055", -- fa58
		x"6100b030", -- fa5c
		x"16bc0003", -- fa60
		x"16bc0084", -- fa64
		x"16bc0002", -- fa68
		x"16bc000b", -- fa6c
		x"4ed016bc", -- fa70
		x"000d6100", -- fa74
		x"ff5018bc", -- fa78
		x"00df16bc", -- fa7c
		x"000b6000", -- fa80
		x"ff446100", -- fa84
		x"fde66100", -- fa88
		x"ff023f00", -- fa8c
		x"3f3c001f", -- fa90
		x"61866100", -- fa94
		x"ff341014", -- fa98
		x"08010003", -- fa9c
		x"6660e148", -- faa0
		x"6100ff26", -- faa4
		x"16bc0083", -- faa8
		x"10143f40", -- faac
		x"000416bc", -- fab0
		x"000d6100", -- fab4
		x"febc803c", -- fab8
		x"00406100", -- fabc
		x"feda6100", -- fac0
		x"ff041880", -- fac4
		x"16bc008a", -- fac8
		x"16bc000b", -- facc
		x"6000fef6", -- fad0
		x"4e560000", -- fad4
		x"6100fd94", -- fad8
		x"3f2e000e", -- fadc
		x"6100feac", -- fae0
		x"3f006100", -- fae4
		x"ff34206e", -- fae8
		x"000a302e", -- faec
		x"00086100", -- faf0
		x"fed85340", -- faf4
		x"6f1610d4", -- faf8
		x"08010003", -- fafc
		x"67f016bc", -- fb00
		x"00836100", -- fb04
		x"ff6a7006", -- fb08
		x"6000fd5a", -- fb0c
		x"16bc0083", -- fb10
		x"10946100", -- fb14
		x"ff5a4e5e", -- fb18
		x"205f508f", -- fb1c
		x"4ed04e56", -- fb20
		x"00006100", -- fb24
		x"fd463f2e", -- fb28
		x"00126100", -- fb2c
		x"fe5e3f00", -- fb30
		x"6100fee6", -- fb34
		x"302e0008", -- fb38
		x"53406d20", -- fb3c
		x"74201212", -- fb40
		x"67fcb202", -- fb44
		x"67100201", -- fb48
		x"002867f2", -- fb4c
		x"08010003", -- fb50
		x"67044a14", -- fb54
		x"60a84a14", -- fb58
		x"51c8ffe4", -- fb5c
		x"202e000a", -- fb60
		x"55806d26", -- fb64
		x"2078fed4", -- fb68
		x"08280005", -- fb6c
		x"000b6650", -- fb70
		x"206e000e", -- fb74
		x"74201212", -- fb78
		x"67fcb202", -- fb7c
		x"663010d4", -- fb80
		x"51c8fff4", -- fb84
		x"42405380", -- fb88
		x"6aec0812", -- fb8c
		x"000567fa", -- fb90
		x"206e000e", -- fb94
		x"202e000a", -- fb98
		x"16bc0083", -- fb9c
		x"119408ff", -- fba0
		x"6100fecc", -- fba4
		x"4e5e205f", -- fba8
		x"defc000c", -- fbac
		x"4ed00201", -- fbb0
		x"002867c2", -- fbb4
		x"08010003", -- fbb8
		x"67c41094", -- fbbc
		x"6000ff40", -- fbc0
		x"41f90050", -- fbc4
		x"000020ae", -- fbc8
		x"000e7200", -- fbcc
		x"74003140", -- fbd0
		x"00043142", -- fbd4
		x"0006137c", -- fbd8
		x"00010003", -- fbdc
		x"40e7007c", -- fbe0
		x"070016bc", -- fbe4
		x"00130829", -- fbe8
		x"00060003", -- fbec
		x"67028212", -- fbf0
		x"16bc0093", -- fbf4
		x"46df0801", -- fbf8
		x"00036606", -- fbfc
		x"05280007", -- fc00
		x"66da1342", -- fc04
		x"00030528", -- fc08
		x"00076706", -- fc0c
		x"4a506000", -- fc10
		x"feee303c", -- fc14
		x"00070c68", -- fc18
		x"ffff0004", -- fc1c
		x"6600fdee", -- fc20
		x"42405380", -- fc24
		x"6ea80801", -- fc28
		x"00056600", -- fc2c
		x"ff646000", -- fc30
		x"ff5a6100", -- fc34
		x"fc3616bc", -- fc38
		x"000c6100", -- fc3c
		x"fd8816bc", -- fc40
		x"008e6100", -- fc44
		x"fd464440", -- fc48
		x"5e404878", -- fc4c
		x"00196100", -- fc50
		x"ae3a0129", -- fc54
		x"001d67fa", -- fc58
		x"16bc000e", -- fc5c
		x"16bc000b", -- fc60
		x"4e754e75", -- fc64
		x"3b40fffe", -- fc68
		x"4e4a45e9", -- fc6c
		x"001747e9", -- fc70
		x"001149e9", -- fc74
		x"00154e75", -- fc78
		x"61f07080", -- fc7c
		x"13400001", -- fc80
		x"13400019", -- fc84
		x"13400019", -- fc88
		x"1340001b", -- fc8c
		x"70010812", -- fc90
		x"000367d0", -- fc94
		x"14bc0040", -- fc98
		x"137c00ff", -- fc9c
		x"001314bc", -- fca0
		x"0000137c", -- fca4
		x"00ff001d", -- fca8
		x"14bc0000", -- fcac
		x"137c0090", -- fcb0
		x"00194878", -- fcb4
		x"00646100", -- fcb8
		x"add2137c", -- fcbc
		x"00a00019", -- fcc0
		x"4e7561a6", -- fcc4
		x"3f3c0010", -- fcc8
		x"61446100", -- fccc
		x"007814bc", -- fcd0
		x"008018bc", -- fcd4
		x"00007004", -- fcd8
		x"6160604c", -- fcdc
		x"4e560000", -- fce0
		x"61883f2e", -- fce4
		x"000e6126", -- fce8
		x"206e000a", -- fcec
		x"302e0008", -- fcf0
		x"61525340", -- fcf4
		x"6f0814bc", -- fcf8
		x"00001898", -- fcfc
		x"60f214bc", -- fd00
		x"00801890", -- fd04
		x"61224e5e", -- fd08
		x"205f508f", -- fd0c
		x"4ed0703f", -- fd10
		x"6128705e", -- fd14
		x"61246116", -- fd18
		x"803c0020", -- fd1c
		x"611c205f", -- fd20
		x"7060805f", -- fd24
		x"2f086012", -- fd28
		x"703f610e", -- fd2c
		x"60162078", -- fd30
		x"fed47000", -- fd34
		x"10280061", -- fd38
		x"4e756108", -- fd3c
		x"14bc0040", -- fd40
		x"18804e75", -- fd44
		x"76016002", -- fd48
		x"76020713", -- fd4c
		x"67024e75", -- fd50
		x"08380001", -- fd54
		x"feda6620", -- fd58
		x"487861a8", -- fd5c
		x"48576100", -- fd60
		x"d9de241f", -- fd64
		x"071366e6", -- fd68
		x"2f024857", -- fd6c
		x"61000200", -- fd70
		x"6af0588f", -- fd74
		x"74006004", -- fd78
		x"343c1af0", -- fd7c
		x"071356ca", -- fd80
		x"fffc66ca", -- fd84
		x"70013f00", -- fd88
		x"6100feee", -- fd8c
		x"301f6000", -- fd90
		x"fed4703f", -- fd94
		x"61a4703e", -- fd98
		x"61a0205f", -- fd9c
		x"7040805f", -- fda0
		x"61987060", -- fda4
		x"805f6192", -- fda8
		x"619a4ed0", -- fdac
		x"705f618a", -- fdb0
		x"60926100", -- fdb4
		x"feb66100", -- fdb8
		x"ff763f00", -- fdbc
		x"3f3c001f", -- fdc0
		x"61d014bc", -- fdc4
		x"008018bc", -- fdc8
		x"00026100", -- fdcc
		x"ff7c1014", -- fdd0
		x"08120006", -- fdd4
		x"6642e148", -- fdd8
		x"6100ff6e", -- fddc
		x"10143f40", -- fde0
		x"0004705e", -- fde4
		x"60c84e56", -- fde8
		x"00006100", -- fdec
		x"fe7e3f2e", -- fdf0
		x"000e6100", -- fdf4
		x"ff3a3f00", -- fdf8
		x"6198206e", -- fdfc
		x"000a302e", -- fe00
		x"000814bc", -- fe04
		x"00801880", -- fe08
		x"6100ff3e", -- fe0c
		x"53406f10", -- fe10
		x"10d40812", -- fe14
		x"000667f0", -- fe18
		x"61927006", -- fe1c
		x"6000fe46", -- fe20
		x"10946188", -- fe24
		x"4e5e205f", -- fe28
		x"508f4ed0", -- fe2c
		x"4e560000", -- fe30
		x"6100fe38", -- fe34
		x"3f2e0012", -- fe38
		x"6100fef4", -- fe3c
		x"3f006100", -- fe40
		x"ff52302e", -- fe44
		x"000848c0", -- fe48
		x"d0ae000a", -- fe4c
		x"b0bc0000", -- fe50
		x"01006f0a", -- fe54
		x"14bc00c0", -- fe58
		x"18bc0000", -- fe5c
		x"600614bc", -- fe60
		x"00801880", -- fe64
		x"302e0008", -- fe68
		x"53406d16", -- fe6c
		x"74027601", -- fe70
		x"12130501", -- fe74
		x"66060701", -- fe78
		x"67f6609c", -- fe7c
		x"4a1451c8", -- fe80
		x"fff0202e", -- fe84
		x"000a5380", -- fe88
		x"2078fed4", -- fe8c
		x"08280005", -- fe90
		x"000b6628", -- fe94
		x"206e000e", -- fe98
		x"74027601", -- fe9c
		x"0513670e", -- fea0
		x"10d451c8", -- fea4
		x"fff84240", -- fea8
		x"53806af0", -- feac
		x"60601213", -- feb0
		x"050166ec", -- feb4
		x"070167e4", -- feb8
		x"6000ff5e", -- febc
		x"41f90050", -- fec0
		x"000020ae", -- fec4
		x"000e7400", -- fec8
		x"137c0001", -- fecc
		x"00033140", -- fed0
		x"0004317c", -- fed4
		x"00080006", -- fed8
		x"08130001", -- fedc
		x"66060528", -- fee0
		x"000766f4", -- fee4
		x"76320528", -- fee8
		x"000757cb", -- feec
		x"fffa6706", -- fef0
		x"61526000", -- fef4
		x"ff240c68", -- fef8
		x"ffff0004", -- fefc
		x"67086144", -- ff00
		x"70076000", -- ff04
		x"fe824240", -- ff08
		x"53806cc2", -- ff0c
		x"61360813", -- ff10
		x"00016618", -- ff14
		x"14bc0000", -- ff18
		x"137c0091", -- ff1c
		x"00194878", -- ff20
		x"00646100", -- ff24
		x"ab66137c", -- ff28
		x"00a00019", -- ff2c
		x"08130002", -- ff30
		x"67044a14", -- ff34
		x"60f66100", -- ff38
		x"fe744e5e", -- ff3c
		x"205fdefc", -- ff40
		x"000c4ed0", -- ff44
		x"4a501342", -- ff48
		x"00034e75", -- ff4c
		x"6100fd1c", -- ff50
		x"6100fdf2", -- ff54
		x"6100fdd8", -- ff58
		x"44405e40", -- ff5c
		x"011467fc", -- ff60
		x"4e754ef9", -- ff64
		x"0000452e", -- ff68
		x"4ef90000", -- ff6c
		x"44d84ef9", -- ff70
		x"0000523e", -- ff74
		x"e75838a1", -- ff78
		x"ffffffff", -- ff7c
		x"15000000", -- ff80
		x"0c001a00", -- ff84
		x"00000c00", -- ff88
		x"05000000", -- ff8c
		x"00001100", -- ff90
		x"00000000", -- ff94
		x"1b000000", -- ff98
		x"01000100", -- ff9c
		x"00000000", -- ffa0
		x"0a010000", -- ffa4
		x"00000801", -- ffa8
		x"00000000", -- ffac
		x"00000000", -- ffb0
		x"00000000", -- ffb4
		x"00000000", -- ffb8
		x"00001200", -- ffbc
		x"0000ff00", -- ffc0
		x"25000000", -- ffc4
		x"00000000", -- ffc8
		x"00002800", -- ffcc
		x"00000000", -- ffd0
		x"00000000", -- ffd4
		x"2a000000", -- ffd8
		x"00000000", -- ffdc
		x"00000300", -- ffe0
		x"00001600", -- ffe4
		x"00002101", -- ffe8
		x"14033312", -- ffec
		x"20151510", -- fff0
		x"150f1515", -- fff4
		x"03151521", -- fff8
		x"00151515", -- fffc
		x"13101014", -- 10000
		x"14041515", -- 10004
		x"15150404", -- 10008
		x"00004e56", -- 1000c
		x"fff42d6e", -- 10010
		x"000cfff8", -- 10014
		x"42aefffc", -- 10018
		x"52aefffc", -- 1001c
		x"206efff8", -- 10020
		x"421052ae", -- 10024
		x"fff80cae", -- 10028
		x"000000b6", -- 1002c
		x"fffc6de8", -- 10030
		x"206e000c", -- 10034
		x"41e80004", -- 10038
		x"2d48fff4", -- 1003c
		x"206efff4", -- 10040
		x"7000102e", -- 10044
		x"000a3080", -- 10048
		x"7000102e", -- 1004c
		x"000b3140", -- 10050
		x"00027000", -- 10054
		x"102e0009", -- 10058
		x"31400004", -- 1005c
		x"42680006", -- 10060
		x"42280008", -- 10064
		x"117c0001", -- 10068
		x"00094228", -- 1006c
		x"00364268", -- 10070
		x"007e4e5e", -- 10074
		x"205f504f", -- 10078
		x"4ed00000", -- 1007c
		x"4e56ffc8", -- 10080
		x"4cba0700", -- 10084
		x"ff5a48ae", -- 10088
		x"0700fffa", -- 1008c
		x"206e0008", -- 10090
		x"022e001f", -- 10094
		x"fffb3028", -- 10098
		x"0008eb88", -- 1009c
		x"812efffb", -- 100a0
		x"206e0008", -- 100a4
		x"2d68000e", -- 100a8
		x"ffc8206e", -- 100ac
		x"00083028", -- 100b0
		x"001248c0", -- 100b4
		x"2d40ffcc", -- 100b8
		x"206e0008", -- 100bc
		x"4ca81e00", -- 100c0
		x"001448ae", -- 100c4
		x"1e00ffd0", -- 100c8
		x"1d68001c", -- 100cc
		x"ffd8206e", -- 100d0
		x"00084ca8", -- 100d4
		x"1e00001e", -- 100d8
		x"48ae1e00", -- 100dc
		x"ffda1d68", -- 100e0
		x"0026ffe2", -- 100e4
		x"206e0008", -- 100e8
		x"43eefffa", -- 100ec
		x"2149000e", -- 100f0
		x"206e0008", -- 100f4
		x"317c0006", -- 100f8
		x"0012206e", -- 100fc
		x"000843ee", -- 10100
		x"ffe42149", -- 10104
		x"0014206e", -- 10108
		x"0008217c", -- 1010c
		x"00000016", -- 10110
		x"0018206e", -- 10114
		x"00084228", -- 10118
		x"001c206e", -- 1011c
		x"000842a8", -- 10120
		x"001e206e", -- 10124
		x"000842a8", -- 10128
		x"0022206e", -- 1012c
		x"00084228", -- 10130
		x"00262f2e", -- 10134
		x"00084eb9", -- 10138
		x"000101d6", -- 1013c
		x"206e0008", -- 10140
		x"216effc8", -- 10144
		x"000e206e", -- 10148
		x"0008316e", -- 1014c
		x"ffce0012", -- 10150
		x"206e0008", -- 10154
		x"4cae1e00", -- 10158
		x"ffd048a8", -- 1015c
		x"1e000014", -- 10160
		x"116effd8", -- 10164
		x"001c206e", -- 10168
		x"00084cae", -- 1016c
		x"1e00ffda", -- 10170
		x"48a81e00", -- 10174
		x"001e116e", -- 10178
		x"ffe20026", -- 1017c
		x"206e0008", -- 10180
		x"4a506600", -- 10184
		x"0040102e", -- 10188
		x"ffe4e888", -- 1018c
		x"02800000", -- 10190
		x"00077207", -- 10194
		x"b2806600", -- 10198
		x"0022102e", -- 1019c
		x"ffe40280", -- 101a0
		x"0000000f", -- 101a4
		x"66000014", -- 101a8
		x"102effe6", -- 101ac
		x"02800000", -- 101b0
		x"000f3d40", -- 101b4
		x"000c6000", -- 101b8
		x"00083d7c", -- 101bc
		x"0012000c", -- 101c0
		x"60000008", -- 101c4
		x"3d7c0012", -- 101c8
		x"000c4e5e", -- 101cc
		x"2e9f4e75", -- 101d0
		x"00004e56", -- 101d4
		x"fff642ae", -- 101d8
		x"fffa206e", -- 101dc
		x"000841e8", -- 101e0
		x"00042d48", -- 101e4
		x"fff6206e", -- 101e8
		x"00084268", -- 101ec
		x"0002206e", -- 101f0
		x"00084250", -- 101f4
		x"206efff6", -- 101f8
		x"42680030", -- 101fc
		x"4268002e", -- 10200
		x"42a80032", -- 10204
		x"226e0008", -- 10208
		x"48690004", -- 1020c
		x"4eb90001", -- 10210
		x"474c206e", -- 10214
		x"fff64a68", -- 10218
		x"00306700", -- 1021c
		x"001a3028", -- 10220
		x"0030226e", -- 10224
		x"00087200", -- 10228
		x"45fafdce", -- 1022c
		x"12320000", -- 10230
		x"32816000", -- 10234
		x"00cc206e", -- 10238
		x"fff64a68", -- 1023c
		x"002e6700", -- 10240
		x"00c01d68", -- 10244
		x"002ffffe", -- 10248
		x"102efffe", -- 1024c
		x"e2880280", -- 10250
		x"0000000f", -- 10254
		x"670000aa", -- 10258
		x"102efffe", -- 1025c
		x"e2880280", -- 10260
		x"0000000f", -- 10264
		x"7201b280", -- 10268
		x"66000032", -- 1026c
		x"2268000a", -- 10270
		x"7003b051", -- 10274
		x"67000018", -- 10278
		x"558f2f2e", -- 1027c
		x"00084eba", -- 10280
		x"fdfc206e", -- 10284
		x"0008315f", -- 10288
		x"00026000", -- 1028c
		x"000c206e", -- 10290
		x"0008317c", -- 10294
		x"00120002", -- 10298
		x"6000002e", -- 1029c
		x"102efffe", -- 102a0
		x"e2880280", -- 102a4
		x"0000000f", -- 102a8
		x"7204b280", -- 102ac
		x"66000010", -- 102b0
		x"206e0008", -- 102b4
		x"317c0013", -- 102b8
		x"00026000", -- 102bc
		x"000c206e", -- 102c0
		x"0008317c", -- 102c4
		x"00110002", -- 102c8
		x"206e0008", -- 102cc
		x"700bb068", -- 102d0
		x"00026600", -- 102d4
		x"00147001", -- 102d8
		x"b0aefffa", -- 102dc
		x"6f00000a", -- 102e0
		x"52aefffa", -- 102e4
		x"6000fef4", -- 102e8
		x"206e0008", -- 102ec
		x"30280002", -- 102f0
		x"206e0008", -- 102f4
		x"720043fa", -- 102f8
		x"fcec1231", -- 102fc
		x"00003081", -- 10300
		x"4e5e2e9f", -- 10304
		x"4e750000", -- 10308
		x"4e56fff4", -- 1030c
		x"426efff4", -- 10310
		x"526efff4", -- 10314
		x"4cba1f00", -- 10318
		x"fcb248ae", -- 1031c
		x"1f00fff6", -- 10320
		x"206e0018", -- 10324
		x"022e001f", -- 10328
		x"fff73028", -- 1032c
		x"0008eb88", -- 10330
		x"812efff7", -- 10334
		x"2d6e0014", -- 10338
		x"fff8202e", -- 1033c
		x"00106c06", -- 10340
		x"d0bc0000", -- 10344
		x"00ffe080", -- 10348
		x"1d40fffd", -- 1034c
		x"202e0010", -- 10350
		x"02800000", -- 10354
		x"00ff1d40", -- 10358
		x"fffe206e", -- 1035c
		x"001843ee", -- 10360
		x"fff62149", -- 10364
		x"000e206e", -- 10368
		x"0018317c", -- 1036c
		x"000a0012", -- 10370
		x"206e0018", -- 10374
		x"216e0008", -- 10378
		x"00142f2e", -- 1037c
		x"000c2f2e", -- 10380
		x"00104eb9", -- 10384
		x"000081b0", -- 10388
		x"206e0018", -- 1038c
		x"215f0018", -- 10390
		x"206e0018", -- 10394
		x"4a680082", -- 10398
		x"57c0206e", -- 1039c
		x"00180200", -- 103a0
		x"00011140", -- 103a4
		x"001c206e", -- 103a8
		x"001842a8", -- 103ac
		x"001e206e", -- 103b0
		x"001842a8", -- 103b4
		x"0022206e", -- 103b8
		x"00184228", -- 103bc
		x"00262f2e", -- 103c0
		x"00184eba", -- 103c4
		x"fe0e206e", -- 103c8
		x"00184a50", -- 103cc
		x"57c06700", -- 103d0
		x"00127002", -- 103d4
		x"b06efff4", -- 103d8
		x"5dc06d00", -- 103dc
		x"00066000", -- 103e0
		x"ff304e5e", -- 103e4
		x"205fdefc", -- 103e8
		x"00144ed0", -- 103ec
		x"00004e56", -- 103f0
		x"ffee426e", -- 103f4
		x"fff03d7c", -- 103f8
		x"0001ffee", -- 103fc
		x"526efff0", -- 10400
		x"7001b06e", -- 10404
		x"ffee6600", -- 10408
		x"00124cba", -- 1040c
		x"0700fb8c", -- 10410
		x"48ae0700", -- 10414
		x"fff26000", -- 10418
		x"00287002", -- 1041c
		x"b06effee", -- 10420
		x"66000012", -- 10424
		x"4cba1f03", -- 10428
		x"fb8448ae", -- 1042c
		x"1f03fff2", -- 10430
		x"6000000e", -- 10434
		x"4cba0700", -- 10438
		x"fb5c48ae", -- 1043c
		x"0700fff2", -- 10440
		x"206e0008", -- 10444
		x"022e001f", -- 10448
		x"fff33028", -- 1044c
		x"0008eb88", -- 10450
		x"812efff3", -- 10454
		x"206e0008", -- 10458
		x"117c0001", -- 1045c
		x"000d206e", -- 10460
		x"000843ee", -- 10464
		x"fff22149", -- 10468
		x"000e206e", -- 1046c
		x"0008317c", -- 10470
		x"00060012", -- 10474
		x"206e0008", -- 10478
		x"42a80014", -- 1047c
		x"206e0008", -- 10480
		x"42a80018", -- 10484
		x"206e0008", -- 10488
		x"4228001c", -- 1048c
		x"206e0008", -- 10490
		x"42a8001e", -- 10494
		x"206e0008", -- 10498
		x"42a80022", -- 1049c
		x"206e0008", -- 104a0
		x"42280026", -- 104a4
		x"2f2e0008", -- 104a8
		x"4ebafd28", -- 104ac
		x"302effee", -- 104b0
		x"5340e340", -- 104b4
		x"323b0006", -- 104b8
		x"4efb1002", -- 104bc
		x"00060028", -- 104c0
		x"007e206e", -- 104c4
		x"00084a50", -- 104c8
		x"6600000a", -- 104cc
		x"426effee", -- 104d0
		x"6000000e", -- 104d4
		x"3d7c0002", -- 104d8
		x"ffee3d7c", -- 104dc
		x"0001fff0", -- 104e0
		x"60000078", -- 104e4
		x"206e0008", -- 104e8
		x"4a506600", -- 104ec
		x"00123d7c", -- 104f0
		x"0001ffee", -- 104f4
		x"3d7c0001", -- 104f8
		x"fff06000", -- 104fc
		x"003a206e", -- 10500
		x"00087002", -- 10504
		x"b0680002", -- 10508
		x"6600002c", -- 1050c
		x"206e0008", -- 10510
		x"7013b068", -- 10514
		x"00026600", -- 10518
		x"00122f3c", -- 1051c
		x"000f4240", -- 10520
		x"4eb90001", -- 10524
		x"4b106000", -- 10528
		x"000e3d7c", -- 1052c
		x"0003ffee", -- 10530
		x"3d7c0001", -- 10534
		x"fff06000", -- 10538
		x"0022206e", -- 1053c
		x"00084a50", -- 10540
		x"66000012", -- 10544
		x"3d7c0001", -- 10548
		x"ffee3d7c", -- 1054c
		x"0001fff0", -- 10550
		x"60000008", -- 10554
		x"3d7c0002", -- 10558
		x"ffee4a6e", -- 1055c
		x"ffee57c0", -- 10560
		x"67000012", -- 10564
		x"7002b06e", -- 10568
		x"fff05dc0", -- 1056c
		x"6d000006", -- 10570
		x"6000fe8a", -- 10574
		x"4e5e2e9f", -- 10578
		x"4e750000", -- 1057c
		x"4e56fffa", -- 10580
		x"4cba0700", -- 10584
		x"fa0a48ae", -- 10588
		x"0700fffa", -- 1058c
		x"206e000c", -- 10590
		x"022e001f", -- 10594
		x"fffb3028", -- 10598
		x"0008eb88", -- 1059c
		x"812efffb", -- 105a0
		x"206e000c", -- 105a4
		x"117c0001", -- 105a8
		x"000d02ae", -- 105ac
		x"000000ff", -- 105b0
		x"fffc202e", -- 105b4
		x"0008e188", -- 105b8
		x"81aefffc", -- 105bc
		x"206e000c", -- 105c0
		x"43eefffa", -- 105c4
		x"2149000e", -- 105c8
		x"206e000c", -- 105cc
		x"317c0006", -- 105d0
		x"0012206e", -- 105d4
		x"000c42a8", -- 105d8
		x"0014206e", -- 105dc
		x"000c42a8", -- 105e0
		x"0018206e", -- 105e4
		x"000c4228", -- 105e8
		x"001c206e", -- 105ec
		x"000c42a8", -- 105f0
		x"001e206e", -- 105f4
		x"000c42a8", -- 105f8
		x"0022206e", -- 105fc
		x"000c4228", -- 10600
		x"00262f2e", -- 10604
		x"000c4eba", -- 10608
		x"fbca4e5e", -- 1060c
		x"205f504f", -- 10610
		x"4ed00000", -- 10614
		x"4e56fff8", -- 10618
		x"426efff8", -- 1061c
		x"526efff8", -- 10620
		x"4cba0700", -- 10624
		x"f98248ae", -- 10628
		x"0700fffa", -- 1062c
		x"206e0014", -- 10630
		x"022e001f", -- 10634
		x"fffb3028", -- 10638
		x"0008eb88", -- 1063c
		x"812efffb", -- 10640
		x"02ae0000", -- 10644
		x"00fffffc", -- 10648
		x"202e0010", -- 1064c
		x"e18881ae", -- 10650
		x"fffc206e", -- 10654
		x"0014117c", -- 10658
		x"0001000d", -- 1065c
		x"206e0014", -- 10660
		x"43eefffa", -- 10664
		x"2149000e", -- 10668
		x"206e0014", -- 1066c
		x"317c0006", -- 10670
		x"0012206e", -- 10674
		x"0014216e", -- 10678
		x"00080014", -- 1067c
		x"2f2e000c", -- 10680
		x"2f2e0010", -- 10684
		x"4eb90000", -- 10688
		x"81b0206e", -- 1068c
		x"0014215f", -- 10690
		x"0018206e", -- 10694
		x"00144a68", -- 10698
		x"008257c0", -- 1069c
		x"206e0014", -- 106a0
		x"02000001", -- 106a4
		x"1140001c", -- 106a8
		x"206e0014", -- 106ac
		x"42a8001e", -- 106b0
		x"206e0014", -- 106b4
		x"42a80022", -- 106b8
		x"206e0014", -- 106bc
		x"42280026", -- 106c0
		x"2f2e0014", -- 106c4
		x"4ebafb0c", -- 106c8
		x"206e0014", -- 106cc
		x"4a5057c0", -- 106d0
		x"67000012", -- 106d4
		x"7002b06e", -- 106d8
		x"fff85dc0", -- 106dc
		x"6d000006", -- 106e0
		x"6000ff3a", -- 106e4
		x"4e5e205f", -- 106e8
		x"defc0010", -- 106ec
		x"4ed00000", -- 106f0
		x"4e56fffa", -- 106f4
		x"4cba0700", -- 106f8
		x"f88a48ae", -- 106fc
		x"0700fffa", -- 10700
		x"206e000c", -- 10704
		x"022e001f", -- 10708
		x"fffb3028", -- 1070c
		x"0008eb88", -- 10710
		x"812efffb", -- 10714
		x"1d7cff0c", -- 10718
		x"fffe206e", -- 1071c
		x"000c117c", -- 10720
		x"0001000d", -- 10724
		x"206e000c", -- 10728
		x"43eefffa", -- 1072c
		x"2149000e", -- 10730
		x"206e000c", -- 10734
		x"317c0006", -- 10738
		x"0012206e", -- 1073c
		x"000c216e", -- 10740
		x"00080014", -- 10744
		x"206e000c", -- 10748
		x"217c0000", -- 1074c
		x"000c0018", -- 10750
		x"206e000c", -- 10754
		x"117c0001", -- 10758
		x"001c206e", -- 1075c
		x"000c42a8", -- 10760
		x"001e206e", -- 10764
		x"000c42a8", -- 10768
		x"0022206e", -- 1076c
		x"000c4228", -- 10770
		x"00262f2e", -- 10774
		x"000c4eba", -- 10778
		x"fa5a4e5e", -- 1077c
		x"205f504f", -- 10780
		x"4ed00000", -- 10784
		x"4e56fffa", -- 10788
		x"4cba0700", -- 1078c
		x"f7f048ae", -- 10790
		x"0700fffa", -- 10794
		x"206e000c", -- 10798
		x"022e001f", -- 1079c
		x"fffb3028", -- 107a0
		x"0008eb88", -- 107a4
		x"812efffb", -- 107a8
		x"1d7cff0c", -- 107ac
		x"fffe206e", -- 107b0
		x"000c117c", -- 107b4
		x"0001000d", -- 107b8
		x"206e000c", -- 107bc
		x"43eefffa", -- 107c0
		x"2149000e", -- 107c4
		x"206e000c", -- 107c8
		x"317c0006", -- 107cc
		x"0012206e", -- 107d0
		x"000c42a8", -- 107d4
		x"0014206e", -- 107d8
		x"000c42a8", -- 107dc
		x"0018206e", -- 107e0
		x"000c4228", -- 107e4
		x"001c206e", -- 107e8
		x"000c216e", -- 107ec
		x"0008001e", -- 107f0
		x"206e000c", -- 107f4
		x"217c0000", -- 107f8
		x"000c0022", -- 107fc
		x"206e000c", -- 10800
		x"117c0001", -- 10804
		x"00262f2e", -- 10808
		x"000c4eba", -- 1080c
		x"f9c64e5e", -- 10810
		x"205f504f", -- 10814
		x"4ed00001", -- 10818
		x"4e56fff2", -- 1081c
		x"206e0008", -- 10820
		x"2d68fffc", -- 10824
		x"fff242ae", -- 10828
		x"fffc52ae", -- 1082c
		x"fffc206e", -- 10830
		x"fff2202e", -- 10834
		x"fffcd080", -- 10838
		x"43e80108", -- 1083c
		x"42710800", -- 10840
		x"0cae0000", -- 10844
		x"0003fffc", -- 10848
		x"6de0206e", -- 1084c
		x"fff22d68", -- 10850
		x"0082fff8", -- 10854
		x"226e0008", -- 10858
		x"2f290008", -- 1085c
		x"2f2efff8", -- 10860
		x"4eb90000", -- 10864
		x"81a8206e", -- 10868
		x"0008215f", -- 1086c
		x"fff82f28", -- 10870
		x"00082f2e", -- 10874
		x"fff84eb9", -- 10878
		x"000081ac", -- 1087c
		x"2d5ffffc", -- 10880
		x"4aaefffc", -- 10884
		x"66000056", -- 10888
		x"206e0008", -- 1088c
		x"2028000c", -- 10890
		x"b0aefff8", -- 10894
		x"6d000046", -- 10898
		x"206e0008", -- 1089c
		x"2f28000c", -- 108a0
		x"2f2efff8", -- 108a4
		x"4eb90000", -- 108a8
		x"81a8206e", -- 108ac
		x"0008215f", -- 108b0
		x"fff42f2e", -- 108b4
		x"fff82f28", -- 108b8
		x"fff44eb9", -- 108bc
		x"000081b0", -- 108c0
		x"206e0008", -- 108c4
		x"215ffff0", -- 108c8
		x"2028fff0", -- 108cc
		x"91a8000c", -- 108d0
		x"2028fff0", -- 108d4
		x"d1a80008", -- 108d8
		x"600000bc", -- 108dc
		x"3d7c0001", -- 108e0
		x"fff6206e", -- 108e4
		x"0008217c", -- 108e8
		x"00000001", -- 108ec
		x"fff44aae", -- 108f0
		x"fffc6f00", -- 108f4
		x"002a202e", -- 108f8
		x"fffc4480", -- 108fc
		x"226efff2", -- 10900
		x"322efff6", -- 10904
		x"48c1d281", -- 10908
		x"45e90108", -- 1090c
		x"35801800", -- 10910
		x"202efffc", -- 10914
		x"91aefff8", -- 10918
		x"3d7c0002", -- 1091c
		x"fff6206e", -- 10920
		x"0008202e", -- 10924
		x"fff8b0a8", -- 10928
		x"000c6d00", -- 1092c
		x"000c2168", -- 10930
		x"000cfff0", -- 10934
		x"6000000c", -- 10938
		x"206e0008", -- 1093c
		x"216efff8", -- 10940
		x"fff0206e", -- 10944
		x"0008226e", -- 10948
		x"fff2302e", -- 1094c
		x"fff648c0", -- 10950
		x"d08045e9", -- 10954
		x"010835a8", -- 10958
		x"fff20800", -- 1095c
		x"526efff6", -- 10960
		x"2028fff0", -- 10964
		x"91a8000c", -- 10968
		x"2028fff0", -- 1096c
		x"d1a80008", -- 10970
		x"2028fff0", -- 10974
		x"91aefff8", -- 10978
		x"4aaefff8", -- 1097c
		x"6f000018", -- 10980
		x"202efff8", -- 10984
		x"4480322e", -- 10988
		x"fff648c1", -- 1098c
		x"d28145e9", -- 10990
		x"01083580", -- 10994
		x"18004e5e", -- 10998
		x"2e9f4e75", -- 1099c
		x"00004e56", -- 109a0
		x"ffec558f", -- 109a4
		x"4eb90000", -- 109a8
		x"aa18301f", -- 109ac
		x"0240001f", -- 109b0
		x"7207b240", -- 109b4
		x"6700000a", -- 109b8
		x"3b7c0001", -- 109bc
		x"fffe4e4a", -- 109c0
		x"2079ffff", -- 109c4
		x"fed42d68", -- 109c8
		x"0010fffc", -- 109cc
		x"202e0008", -- 109d0
		x"e1802d40", -- 109d4
		x"00084aae", -- 109d8
		x"000c6f00", -- 109dc
		x"00e42d6e", -- 109e0
		x"fffcffec", -- 109e4
		x"206effec", -- 109e8
		x"48680088", -- 109ec
		x"2279ffff", -- 109f0
		x"fed42f29", -- 109f4
		x"005e4eba", -- 109f8
		x"f6122f0e", -- 109fc
		x"4ebafe1a", -- 10a00
		x"2079ffff", -- 10a04
		x"fed41028", -- 10a08
		x"005e0280", -- 10a0c
		x"0000001f", -- 10a10
		x"720fb280", -- 10a14
		x"66000050", -- 10a18
		x"206effec", -- 10a1c
		x"202efff8", -- 10a20
		x"b0a8007e", -- 10a24
		x"67000014", -- 10a28
		x"48680088", -- 10a2c
		x"202efff8", -- 10a30
		x"90a8007e", -- 10a34
		x"2f004eba", -- 10a38
		x"fb44206e", -- 10a3c
		x"ffec4868", -- 10a40
		x"00882f2e", -- 10a44
		x"fff42f28", -- 10a48
		x"00822f2e", -- 10a4c
		x"00104eba", -- 10a50
		x"fbc4202e", -- 10a54
		x"fff8d0ae", -- 10a58
		x"fff4206e", -- 10a5c
		x"ffec2140", -- 10a60
		x"007e6000", -- 10a64
		x"003c202e", -- 10a68
		x"fff8d0ae", -- 10a6c
		x"fff45380", -- 10a70
		x"206effec", -- 10a74
		x"b0a8007e", -- 10a78
		x"6f00000a", -- 10a7c
		x"3b7c0004", -- 10a80
		x"fffe4e4a", -- 10a84
		x"206effec", -- 10a88
		x"48680088", -- 10a8c
		x"2f2efff8", -- 10a90
		x"2f2efff4", -- 10a94
		x"2f280082", -- 10a98
		x"2f2e0010", -- 10a9c
		x"4ebaf86a", -- 10aa0
		x"206effec", -- 10aa4
		x"4a680088", -- 10aa8
		x"6700000a", -- 10aac
		x"3b7c0004", -- 10ab0
		x"fffe4e4a", -- 10ab4
		x"202efff0", -- 10ab8
		x"d1ae0010", -- 10abc
		x"6000ff18", -- 10ac0
		x"4e5e205f", -- 10ac4
		x"defc000c", -- 10ac8
		x"4ed00000", -- 10acc
		x"4e56ffde", -- 10ad0
		x"2d6e0008", -- 10ad4
		x"fff62f2d", -- 10ad8
		x"fff62f0e", -- 10adc
		x"487a01d6", -- 10ae0
		x"2b4ffff6", -- 10ae4
		x"2079ffff", -- 10ae8
		x"fed47000", -- 10aec
		x"10280060", -- 10af0
		x"3f004eb9", -- 10af4
		x"00011902", -- 10af8
		x"4cba0700", -- 10afc
		x"f4be48ae", -- 10b00
		x"0700fffa", -- 10b04
		x"2079ffff", -- 10b08
		x"fed41028", -- 10b0c
		x"005f022e", -- 10b10
		x"001ffffb", -- 10b14
		x"eb080200", -- 10b18
		x"00e0812e", -- 10b1c
		x"fffb1d7c", -- 10b20
		x"fffffffe", -- 10b24
		x"2079ffff", -- 10b28
		x"fed42d68", -- 10b2c
		x"0010ffde", -- 10b30
		x"206effde", -- 10b34
		x"48680088", -- 10b38
		x"2279ffff", -- 10b3c
		x"fed42f29", -- 10b40
		x"005e4eba", -- 10b44
		x"f4c6206e", -- 10b48
		x"ffde43ee", -- 10b4c
		x"fffa2149", -- 10b50
		x"0096317c", -- 10b54
		x"0006009a", -- 10b58
		x"216efff6", -- 10b5c
		x"009c7000", -- 10b60
		x"102efffe", -- 10b64
		x"214000a0", -- 10b68
		x"422800a4", -- 10b6c
		x"42a800a6", -- 10b70
		x"42a800aa", -- 10b74
		x"422800ae", -- 10b78
		x"48680088", -- 10b7c
		x"4ebaf654", -- 10b80
		x"206effde", -- 10b84
		x"4a680088", -- 10b88
		x"66000108", -- 10b8c
		x"226efff6", -- 10b90
		x"08290007", -- 10b94
		x"000156c0", -- 10b98
		x"44001d40", -- 10b9c
		x"ffe3226e", -- 10ba0
		x"fff67000", -- 10ba4
		x"10290004", -- 10ba8
		x"0c4000fa", -- 10bac
		x"6f00000c", -- 10bb0
		x"226efff6", -- 10bb4
		x"137cfffa", -- 10bb8
		x"000441fa", -- 10bbc
		x"01261018", -- 10bc0
		x"43eeffe4", -- 10bc4
		x"12c012d8", -- 10bc8
		x"530062fa", -- 10bcc
		x"1f3cff10", -- 10bd0
		x"486effe4", -- 10bd4
		x"2f3c0000", -- 10bd8
		x"0001206e", -- 10bdc
		x"fff61f3c", -- 10be0
		x"fffa4868", -- 10be4
		x"00042f3c", -- 10be8
		x"0000000c", -- 10bec
		x"2f3c0000", -- 10bf0
		x"00104eb9", -- 10bf4
		x"000081fe", -- 10bf8
		x"1f3c00ff", -- 10bfc
		x"2f2e0008", -- 10c00
		x"2f3c0000", -- 10c04
		x"0001206e", -- 10c08
		x"fff61f3c", -- 10c0c
		x"fffa4868", -- 10c10
		x"00042f3c", -- 10c14
		x"00000004", -- 10c18
		x"2f3c0000", -- 10c1c
		x"00084eb9", -- 10c20
		x"000081fe", -- 10c24
		x"1f3c00ff", -- 10c28
		x"2f2e0008", -- 10c2c
		x"4eb90001", -- 10c30
		x"4bb8206e", -- 10c34
		x"00087000", -- 10c38
		x"10105240", -- 10c3c
		x"206e0008", -- 10c40
		x"1080206e", -- 10c44
		x"0008226e", -- 10c48
		x"00087000", -- 10c4c
		x"101111bc", -- 10c50
		x"00200000", -- 10c54
		x"1f3c00ff", -- 10c58
		x"2f2e0008", -- 10c5c
		x"486effe4", -- 10c60
		x"4eb90000", -- 10c64
		x"81cc1f3c", -- 10c68
		x"00ff2f2e", -- 10c6c
		x"00084eb9", -- 10c70
		x"00014bb8", -- 10c74
		x"4a2effe3", -- 10c78
		x"67000014", -- 10c7c
		x"1f3c00ff", -- 10c80
		x"2f2e0008", -- 10c84
		x"487a005e", -- 10c88
		x"4eb90000", -- 10c8c
		x"81cc6000", -- 10c90
		x"001641fa", -- 10c94
		x"00561018", -- 10c98
		x"246e0008", -- 10c9c
		x"43d212c0", -- 10ca0
		x"12d85300", -- 10ca4
		x"62fa2b6f", -- 10ca8
		x"0008fff6", -- 10cac
		x"defc000c", -- 10cb0
		x"4efa002a", -- 10cb4
		x"2c5f2b5f", -- 10cb8
		x"fff641fa", -- 10cbc
		x"00361018", -- 10cc0
		x"246e0008", -- 10cc4
		x"43d212c0", -- 10cc8
		x"12d85300", -- 10ccc
		x"62fa7030", -- 10cd0
		x"d06dfffe", -- 10cd4
		x"206e0008", -- 10cd8
		x"1140000d", -- 10cdc
		x"4e5e2e9f", -- 10ce0
		x"4e750000", -- 10ce4
		x"05205245", -- 10ce8
		x"4d560775", -- 10cec
		x"6e6b6e6f", -- 10cf0
		x"776e0d75", -- 10cf4
		x"6e6b6e6f", -- 10cf8
		x"776e2c20", -- 10cfc
		x"65633d20", -- 10d00
		x"00004e56", -- 10d04
		x"ffea2079", -- 10d08
		x"fffffed4", -- 10d0c
		x"2d680010", -- 10d10
		x"fff02d6e", -- 10d14
		x"fff0ffea", -- 10d18
		x"206effea", -- 10d1c
		x"217cffff", -- 10d20
		x"ffff0082", -- 10d24
		x"42a8007e", -- 10d28
		x"558f4eb9", -- 10d2c
		x"0001120c", -- 10d30
		x"206effea", -- 10d34
		x"315f0086", -- 10d38
		x"558f3f3c", -- 10d3c
		x"00073f28", -- 10d40
		x"00864eb9", -- 10d44
		x"00011048", -- 10d48
		x"4a1f6600", -- 10d4c
		x"000a3b7c", -- 10d50
		x"0001fffe", -- 10d54
		x"4e4a206e", -- 10d58
		x"ffea4868", -- 10d5c
		x"00882279", -- 10d60
		x"fffffed4", -- 10d64
		x"2f29005e", -- 10d68
		x"4ebaf2a0", -- 10d6c
		x"206effea", -- 10d70
		x"48680088", -- 10d74
		x"4ebaf678", -- 10d78
		x"206effea", -- 10d7c
		x"4a680088", -- 10d80
		x"67000020", -- 10d84
		x"7013b068", -- 10d88
		x"008a6600", -- 10d8c
		x"000e3b7c", -- 10d90
		x"0003fffe", -- 10d94
		x"4e4a6000", -- 10d98
		x"000a3b7c", -- 10d9c
		x"0002fffe", -- 10da0
		x"4e4a426e", -- 10da4
		x"ffee526e", -- 10da8
		x"ffee206e", -- 10dac
		x"ffea4868", -- 10db0
		x"00882279", -- 10db4
		x"fffffed4", -- 10db8
		x"2f29005e", -- 10dbc
		x"4ebaf24c", -- 10dc0
		x"206effea", -- 10dc4
		x"48680088", -- 10dc8
		x"486efff4", -- 10dcc
		x"4ebaf922", -- 10dd0
		x"206effea", -- 10dd4
		x"4a680088", -- 10dd8
		x"660000bc", -- 10ddc
		x"202efffc", -- 10de0
		x"028000ff", -- 10de4
		x"ffff6600", -- 10de8
		x"001402ae", -- 10dec
		x"ff000000", -- 10df0
		x"fffc203c", -- 10df4
		x"00000100", -- 10df8
		x"81aefffc", -- 10dfc
		x"202efffc", -- 10e00
		x"028000ff", -- 10e04
		x"ffff0c80", -- 10e08
		x"00000100", -- 10e0c
		x"6c00000a", -- 10e10
		x"3b7c0001", -- 10e14
		x"fffe4e4a", -- 10e18
		x"558f202e", -- 10e1c
		x"fffc0280", -- 10e20
		x"00ffffff", -- 10e24
		x"2f004eb9", -- 10e28
		x"00014b72", -- 10e2c
		x"4a1f6600", -- 10e30
		x"000a3b7c", -- 10e34
		x"0001fffe", -- 10e38
		x"4e4a206e", -- 10e3c
		x"ffea202e", -- 10e40
		x"fffc0280", -- 10e44
		x"00ffffff", -- 10e48
		x"21400082", -- 10e4c
		x"102efff6", -- 10e50
		x"e8880280", -- 10e54
		x"00000007", -- 10e58
		x"6700003c", -- 10e5c
		x"1d7c0000", -- 10e60
		x"fff41d7c", -- 10e64
		x"0000fff5", -- 10e68
		x"08ae0007", -- 10e6c
		x"fff6022e", -- 10e70
		x"008ffff6", -- 10e74
		x"7000e988", -- 10e78
		x"812efff6", -- 10e7c
		x"02aeff00", -- 10e80
		x"0000fff8", -- 10e84
		x"700081ae", -- 10e88
		x"fff84868", -- 10e8c
		x"0088486e", -- 10e90
		x"fff44eba", -- 10e94
		x"f8f0206e", -- 10e98
		x"ffea4a68", -- 10e9c
		x"008857c0", -- 10ea0
		x"67000012", -- 10ea4
		x"7002b06e", -- 10ea8
		x"ffee5dc0", -- 10eac
		x"6d000006", -- 10eb0
		x"6000fef4", -- 10eb4
		x"206effea", -- 10eb8
		x"4a680088", -- 10ebc
		x"6700000a", -- 10ec0
		x"3b7c0001", -- 10ec4
		x"fffe4e4a", -- 10ec8
		x"4e5e4e75", -- 10ecc
		x"00004e56", -- 10ed0
		x"ffe02079", -- 10ed4
		x"fffffed4", -- 10ed8
		x"2d680010", -- 10edc
		x"ffea2d6e", -- 10ee0
		x"ffeaffe4", -- 10ee4
		x"558f4eb9", -- 10ee8
		x"0001120c", -- 10eec
		x"206effe4", -- 10ef0
		x"315f0086", -- 10ef4
		x"558f3f3c", -- 10ef8
		x"00073f28", -- 10efc
		x"00864eb9", -- 10f00
		x"0001109c", -- 10f04
		x"4a1f6600", -- 10f08
		x"000a3b7c", -- 10f0c
		x"0001fffe", -- 10f10
		x"4e4a4cba", -- 10f14
		x"1f00f0aa", -- 10f18
		x"48ae1f00", -- 10f1c
		x"fff62079", -- 10f20
		x"fffffed4", -- 10f24
		x"1028005f", -- 10f28
		x"022e001f", -- 10f2c
		x"fff7eb08", -- 10f30
		x"020000e0", -- 10f34
		x"812efff7", -- 10f38
		x"426effe8", -- 10f3c
		x"206effe4", -- 10f40
		x"48680088", -- 10f44
		x"2279ffff", -- 10f48
		x"fed42f29", -- 10f4c
		x"005e4eba", -- 10f50
		x"f0ba206e", -- 10f54
		x"ffe443ee", -- 10f58
		x"fff62149", -- 10f5c
		x"0096317c", -- 10f60
		x"000a009a", -- 10f64
		x"43eeffee", -- 10f68
		x"2149009c", -- 10f6c
		x"217c0000", -- 10f70
		x"000800a0", -- 10f74
		x"422800a4", -- 10f78
		x"42a800a6", -- 10f7c
		x"42a800aa", -- 10f80
		x"422800ae", -- 10f84
		x"48680088", -- 10f88
		x"4ebaf248", -- 10f8c
		x"526effe8", -- 10f90
		x"206effe4", -- 10f94
		x"4a680088", -- 10f98
		x"57c06700", -- 10f9c
		x"00107003", -- 10fa0
		x"b06effe8", -- 10fa4
		x"5dc06d00", -- 10fa8
		x"00046090", -- 10fac
		x"206effe4", -- 10fb0
		x"4a680088", -- 10fb4
		x"66000054", -- 10fb8
		x"43e8007e", -- 10fbc
		x"2d49ffe0", -- 10fc0
		x"7020b0ae", -- 10fc4
		x"fff26e00", -- 10fc8
		x"002e0cae", -- 10fcc
		x"00100000", -- 10fd0
		x"fff26e00", -- 10fd4
		x"0022558f", -- 10fd8
		x"2f2efff2", -- 10fdc
		x"4eb90001", -- 10fe0
		x"4b724a1f", -- 10fe4
		x"67000010", -- 10fe8
		x"206effe0", -- 10fec
		x"216efff2", -- 10ff0
		x"00046000", -- 10ff4
		x"000a3b7c", -- 10ff8
		x"0002fffe", -- 10ffc
		x"4e4a206e", -- 11000
		x"ffe020ae", -- 11004
		x"ffee6000", -- 11008
		x"0036206e", -- 1100c
		x"ffe47013", -- 11010
		x"b068008a", -- 11014
		x"57c06700", -- 11018
		x"00127002", -- 1101c
		x"b068008a", -- 11020
		x"57c06700", -- 11024
		x"00066000", -- 11028
		x"000e3b7c", -- 1102c
		x"0003fffe", -- 11030
		x"4e4a6000", -- 11034
		x"000a3b7c", -- 11038
		x"0001fffe", -- 1103c
		x"4e4a4e5e", -- 11040
		x"4e750000", -- 11044
		x"4e56fffe", -- 11048
		x"3d6e0008", -- 1104c
		x"fffe322e", -- 11050
		x"000a0241", -- 11054
		x"001f7407", -- 11058
		x"b44157c1", -- 1105c
		x"10016700", -- 11060
		x"00282079", -- 11064
		x"fffffed4", -- 11068
		x"1228005e", -- 1106c
		x"02810000", -- 11070
		x"001f740f", -- 11074
		x"b48157c1", -- 11078
		x"10016700", -- 1107c
		x"000c7201", -- 11080
		x"b22efffe", -- 11084
		x"57c11001", -- 11088
		x"0200ff01", -- 1108c
		x"1d40000c", -- 11090
		x"4e5e2e9f", -- 11094
		x"4e750000", -- 11098
		x"4e56fffa", -- 1109c
		x"3d6e0008", -- 110a0
		x"fffe322e", -- 110a4
		x"000a0241", -- 110a8
		x"001f7407", -- 110ac
		x"b44157c1", -- 110b0
		x"10016700", -- 110b4
		x"003a2079", -- 110b8
		x"fffffed4", -- 110bc
		x"1228005e", -- 110c0
		x"02810000", -- 110c4
		x"001f740e", -- 110c8
		x"b48157c1", -- 110cc
		x"10016700", -- 110d0
		x"001e7200", -- 110d4
		x"122efffe", -- 110d8
		x"2f01487a", -- 110dc
		x"00202d40", -- 110e0
		x"fffa4eb9", -- 110e4
		x"000081b4", -- 110e8
		x"202efffa", -- 110ec
		x"101f0200", -- 110f0
		x"ff011d40", -- 110f4
		x"000c4e5e", -- 110f8
		x"2e9f4e75", -- 110fc
		x"00028d00", -- 11100
		x"00004e56", -- 11104
		x"fffc2d79", -- 11108
		x"fffffed4", -- 1110c
		x"fffc206e", -- 11110
		x"fffc7000", -- 11114
		x"10280060", -- 11118
		x"3f004eb9", -- 1111c
		x"00011902", -- 11120
		x"4a2e0008", -- 11124
		x"67000018", -- 11128
		x"206efffc", -- 1112c
		x"70001028", -- 11130
		x"00603f00", -- 11134
		x"4eb90001", -- 11138
		x"236a6000", -- 1113c
		x"0014206e", -- 11140
		x"fffc7000", -- 11144
		x"10280060", -- 11148
		x"3f004eb9", -- 1114c
		x"0001227e", -- 11150
		x"4e5e205f", -- 11154
		x"544f4ed0", -- 11158
		x"00004e56", -- 1115c
		x"00004227", -- 11160
		x"4ebaffa0", -- 11164
		x"4e5e4e75", -- 11168
		x"00004e56", -- 1116c
		x"fff82d79", -- 11170
		x"fffffed4", -- 11174
		x"fff82f3c", -- 11178
		x"00010000", -- 1117c
		x"206efff8", -- 11180
		x"70001028", -- 11184
		x"00607260", -- 11188
		x"d24048c1", -- 1118c
		x"2f014eb9", -- 11190
		x"000081b0", -- 11194
		x"2d5ffffc", -- 11198
		x"206efff8", -- 1119c
		x"4a28005f", -- 111a0
		x"54c11001", -- 111a4
		x"67000054", -- 111a8
		x"7207b228", -- 111ac
		x"005f54c1", -- 111b0
		x"10016700", -- 111b4
		x"0046206e", -- 111b8
		x"fff84a28", -- 111bc
		x"006154c1", -- 111c0
		x"10016700", -- 111c4
		x"0036206e", -- 111c8
		x"fff87207", -- 111cc
		x"b2280061", -- 111d0
		x"54c11001", -- 111d4
		x"67000024", -- 111d8
		x"206efffc", -- 111dc
		x"12280007", -- 111e0
		x"02810000", -- 111e4
		x"00077407", -- 111e8
		x"9481206e", -- 111ec
		x"fff87200", -- 111f0
		x"12280061", -- 111f4
		x"b28256c1", -- 111f8
		x"10010200", -- 111fc
		x"00011d40", -- 11200
		x"00084e5e", -- 11204
		x"4e750000", -- 11208
		x"4e56fff0", -- 1120c
		x"3d7cffff", -- 11210
		x"0008558f", -- 11214
		x"4eb90000", -- 11218
		x"aa18301f", -- 1121c
		x"0240001f", -- 11220
		x"7207b240", -- 11224
		x"6700000a", -- 11228
		x"3b7c0001", -- 1122c
		x"fffe4e4a", -- 11230
		x"558f4eba", -- 11234
		x"ff364a1f", -- 11238
		x"670000d4", -- 1123c
		x"2d79ffff", -- 11240
		x"fed4fff4", -- 11244
		x"206efff4", -- 11248
		x"2d680010", -- 1124c
		x"fff07000", -- 11250
		x"10280060", -- 11254
		x"3f004eb9", -- 11258
		x"00011902", -- 1125c
		x"42a74879", -- 11260
		x"0001490e", -- 11264
		x"206efff4", -- 11268
		x"70001028", -- 1126c
		x"00603f00", -- 11270
		x"4eb90001", -- 11274
		x"1a4e206e", -- 11278
		x"fff47000", -- 1127c
		x"10280060", -- 11280
		x"3f004eb9", -- 11284
		x"0001227e", -- 11288
		x"4cba0700", -- 1128c
		x"ed2e48ae", -- 11290
		x"0700fff8", -- 11294
		x"206efff4", -- 11298
		x"1028005f", -- 1129c
		x"022e001f", -- 112a0
		x"fff9eb08", -- 112a4
		x"020000e0", -- 112a8
		x"812efff9", -- 112ac
		x"1d7cff02", -- 112b0
		x"fffc226e", -- 112b4
		x"fff04869", -- 112b8
		x"00882f28", -- 112bc
		x"005e4eba", -- 112c0
		x"ed4a206e", -- 112c4
		x"fff043ee", -- 112c8
		x"fff82149", -- 112cc
		x"0096317c", -- 112d0
		x"0006009a", -- 112d4
		x"43eefffe", -- 112d8
		x"2149009c", -- 112dc
		x"217c0000", -- 112e0
		x"000200a0", -- 112e4
		x"422800a4", -- 112e8
		x"42a800a6", -- 112ec
		x"42a800aa", -- 112f0
		x"422800ae", -- 112f4
		x"48680088", -- 112f8
		x"4ebaeed8", -- 112fc
		x"206efff0", -- 11300
		x"4a680088", -- 11304
		x"66000008", -- 11308
		x"3d6efffe", -- 1130c
		x"00084e5e", -- 11310
		x"4e754e75", -- 11314
		x"30cb27b9", -- 11318
		x"ffffffff", -- 1131c
		x"205f201f", -- 11320
		x"221f225f", -- 11324
		x"42290011", -- 11328
		x"23410016", -- 1132c
		x"23410012", -- 11330
		x"2340001a", -- 11334
		x"4ed0205f", -- 11338
		x"101f225f", -- 1133c
		x"13400011", -- 11340
		x"670c4aa9", -- 11344
		x"00126e00", -- 11348
		x"00064229", -- 1134c
		x"00114ed0", -- 11350
		x"4e56fffc", -- 11354
		x"206e0014", -- 11358
		x"216e0010", -- 1135c
		x"0000216e", -- 11360
		x"000c0004", -- 11364
		x"42a80008", -- 11368
		x"4268000c", -- 1136c
		x"4268000e", -- 11370
		x"42280010", -- 11374
		x"42280011", -- 11378
		x"42a80012", -- 1137c
		x"216e0008", -- 11380
		x"001e42a8", -- 11384
		x"00224e5e", -- 11388
		x"205fdefc", -- 1138c
		x"00104ed0", -- 11390
		x"4e56fffc", -- 11394
		x"2d6e000c", -- 11398
		x"fffc206e", -- 1139c
		x"fffc216e", -- 113a0
		x"00080000", -- 113a4
		x"42a80008", -- 113a8
		x"4268000c", -- 113ac
		x"4268000e", -- 113b0
		x"42280010", -- 113b4
		x"42280011", -- 113b8
		x"21680016", -- 113bc
		x"00124aa8", -- 113c0
		x"00226706", -- 113c4
		x"21680026", -- 113c8
		x"000442a8", -- 113cc
		x"00224e5e", -- 113d0
		x"205f504f", -- 113d4
		x"4ed04e56", -- 113d8
		x"fff4206e", -- 113dc
		x"00082d68", -- 113e0
		x"0008fffc", -- 113e4
		x"226efffc", -- 113e8
		x"2469001a", -- 113ec
		x"20290012", -- 113f0
		x"2f002f3c", -- 113f4
		x"00000006", -- 113f8
		x"2d4afff8", -- 113fc
		x"4eb90000", -- 11400
		x"81b0246e", -- 11404
		x"fff8201f", -- 11408
		x"41f208fa", -- 1140c
		x"2d48fff4", -- 11410
		x"206efff4", -- 11414
		x"30ae000c", -- 11418
		x"30106d52", -- 1141c
		x"b07c0003", -- 11420
		x"6e4ce340", -- 11424
		x"323b0006", -- 11428
		x"4efb1002", -- 1142c
		x"00080024", -- 11430
		x"00140034", -- 11434
		x"226efffc", -- 11438
		x"21690008", -- 1143c
		x"0002602e", -- 11440
		x"206efffc", -- 11444
		x"226efff4", -- 11448
		x"23680004", -- 1144c
		x"0002601e", -- 11450
		x"206e0008", -- 11454
		x"226efff4", -- 11458
		x"2368ffe6", -- 1145c
		x"0002600e", -- 11460
		x"206e0008", -- 11464
		x"226efff4", -- 11468
		x"2368ffee", -- 1146c
		x"0002206e", -- 11470
		x"fffc53a8", -- 11474
		x"00124aa8", -- 11478
		x"00125ec0", -- 1147c
		x"02000001", -- 11480
		x"11400011", -- 11484
		x"4e5e205f", -- 11488
		x"5c4f4ed0", -- 1148c
		x"4e56fffa", -- 11490
		x"122e000c", -- 11494
		x"206e0008", -- 11498
		x"22680008", -- 1149c
		x"4a69000c", -- 114a0
		x"663270fb", -- 114a4
		x"b0416706", -- 114a8
		x"70fdb041", -- 114ac
		x"66263341", -- 114b0
		x"000c70fb", -- 114b4
		x"b0416608", -- 114b8
		x"336dfffe", -- 114bc
		x"000e6006", -- 114c0
		x"3368fff0", -- 114c4
		x"000e2469", -- 114c8
		x"00047000", -- 114cc
		x"30122140", -- 114d0
		x"0008600e", -- 114d4
		x"137c0001", -- 114d8
		x"00104228", -- 114dc
		x"ffff3341", -- 114e0
		x"000c4e5e", -- 114e4
		x"205f5c4f", -- 114e8
		x"4ed04e56", -- 114ec
		x"fff8206e", -- 114f0
		x"00082468", -- 114f4
		x"00082d4a", -- 114f8
		x"fffc2268", -- 114fc
		x"fffa2d49", -- 11500
		x"fff87000", -- 11504
		x"10290001", -- 11508
		x"6d0000b0", -- 1150c
		x"b07c0003", -- 11510
		x"6e0000a8", -- 11514
		x"e340323b", -- 11518
		x"00064efb", -- 1151c
		x"10020008", -- 11520
		x"0008004c", -- 11524
		x"004c7000", -- 11528
		x"10290002", -- 1152c
		x"b0a8ffee", -- 11530
		x"6f142028", -- 11534
		x"ffeed080", -- 11538
		x"72003231", -- 1153c
		x"08042541", -- 11540
		x"00086000", -- 11544
		x"00827201", -- 11548
		x"b2290001", -- 1154c
		x"66145340", -- 11550
		x"48c0d080", -- 11554
		x"72003230", -- 11558
		x"08042541", -- 1155c
		x"00086000", -- 11560
		x"00663f3c", -- 11564
		x"fffd6000", -- 11568
		x"00564287", -- 1156c
		x"70001029", -- 11570
		x"0002b087", -- 11574
		x"6f242007", -- 11578
		x"e5807200", -- 1157c
		x"32310804", -- 11580
		x"b2a8ffee", -- 11584
		x"6610e587", -- 11588
		x"72003231", -- 1158c
		x"78062541", -- 11590
		x"00086000", -- 11594
		x"00325287", -- 11598
		x"60d27203", -- 1159c
		x"b2290001", -- 115a0
		x"66125340", -- 115a4
		x"48c0e580", -- 115a8
		x"72003231", -- 115ac
		x"08062541", -- 115b0
		x"00086012", -- 115b4
		x"3f3cfffd", -- 115b8
		x"60043f3c", -- 115bc
		x"fffe2f2e", -- 115c0
		x"00084eba", -- 115c4
		x"fec84e5e", -- 115c8
		x"2e9f4e75", -- 115cc
		x"4e56ffde", -- 115d0
		x"1d7c0001", -- 115d4
		x"ffff42ae", -- 115d8
		x"fffa206e", -- 115dc
		x"00082d48", -- 115e0
		x"ffe24a28", -- 115e4
		x"0011670a", -- 115e8
		x"3f3c0002", -- 115ec
		x"2f0e4eba", -- 115f0
		x"fde6206e", -- 115f4
		x"ffe24228", -- 115f8
		x"00104aa8", -- 115fc
		x"00086608", -- 11600
		x"217c0000", -- 11604
		x"00020008", -- 11608
		x"206effe2", -- 1160c
		x"20280008", -- 11610
		x"2d680004", -- 11614
		x"fffad1ae", -- 11618
		x"fffa4a28", -- 1161c
		x"00116708", -- 11620
		x"42672f0e", -- 11624
		x"4ebafdb0", -- 11628
		x"206efffa", -- 1162c
		x"2d48ffde", -- 11630
		x"70001028", -- 11634
		x"00006d00", -- 11638
		x"0226b07c", -- 1163c
		x"00046e00", -- 11640
		x"021ee340", -- 11644
		x"323b0006", -- 11648
		x"4efb1002", -- 1164c
		x"000a00fa", -- 11650
		x"01ae01f0", -- 11654
		x"02082f2d", -- 11658
		x"fff62f0e", -- 1165c
		x"487a00d4", -- 11660
		x"2b4ffff6", -- 11664
		x"70001028", -- 11668
		x"00016d44", -- 1166c
		x"b07c0003", -- 11670
		x"6e3ee340", -- 11674
		x"323b0006", -- 11678
		x"4efb1002", -- 1167c
		x"00080008", -- 11680
		x"001c001c", -- 11684
		x"70001028", -- 11688
		x"000248c0", -- 1168c
		x"d08043f0", -- 11690
		x"08042d49", -- 11694
		x"fff66026", -- 11698
		x"206effde", -- 1169c
		x"70001028", -- 116a0
		x"000248c0", -- 116a4
		x"e58043f0", -- 116a8
		x"08042d49", -- 116ac
		x"fff6600e", -- 116b0
		x"3f3cfffe", -- 116b4
		x"2f0e4eba", -- 116b8
		x"fdd46000", -- 116bc
		x"01ac206e", -- 116c0
		x"ffde7000", -- 116c4
		x"10280003", -- 116c8
		x"2d40fff2", -- 116cc
		x"6750206e", -- 116d0
		x"fff62d50", -- 116d4
		x"ffe6206e", -- 116d8
		x"ffe24a28", -- 116dc
		x"0011670e", -- 116e0
		x"3f3c0001", -- 116e4
		x"2f0e4eba", -- 116e8
		x"fcee206e", -- 116ec
		x"ffe22f10", -- 116f0
		x"486effee", -- 116f4
		x"226effe6", -- 116f8
		x"4e91206e", -- 116fc
		x"ffe24a28", -- 11700
		x"0011670a", -- 11704
		x"3f3c0003", -- 11708
		x"2f0e4eba", -- 1170c
		x"fcca4aae", -- 11710
		x"ffee660a", -- 11714
		x"58aefff6", -- 11718
		x"53aefff2", -- 1171c
		x"66b02f0e", -- 11720
		x"4ebafdc8", -- 11724
		x"2b6f0008", -- 11728
		x"fff6defc", -- 1172c
		x"000c6000", -- 11730
		x"01382c5f", -- 11734
		x"2b5ffff6", -- 11738
		x"3f3cfffb", -- 1173c
		x"2f0e4eba", -- 11740
		x"fd4c6000", -- 11744
		x"0124206e", -- 11748
		x"ffe22028", -- 1174c
		x"0022b0a8", -- 11750
		x"001e6c00", -- 11754
		x"009852a8", -- 11758
		x"00222028", -- 1175c
		x"0022e780", -- 11760
		x"21a80004", -- 11764
		x"081e21ae", -- 11768
		x"fffa0822", -- 1176c
		x"226effde", -- 11770
		x"70001029", -- 11774
		x"00016d40", -- 11778
		x"b07c0003", -- 1177c
		x"6e3ae340", -- 11780
		x"323b0006", -- 11784
		x"4efb1002", -- 11788
		x"00080008", -- 1178c
		x"001c001c", -- 11790
		x"70001029", -- 11794
		x"000248c0", -- 11798
		x"d08045f1", -- 1179c
		x"08042d4a", -- 117a0
		x"fff66022", -- 117a4
		x"70001029", -- 117a8
		x"000248c0", -- 117ac
		x"e58045f1", -- 117b0
		x"08042d4a", -- 117b4
		x"fff6600e", -- 117b8
		x"3f3cfffe", -- 117bc
		x"2f0e4eba", -- 117c0
		x"fccc6000", -- 117c4
		x"00a42152", -- 117c8
		x"000442ae", -- 117cc
		x"fffa217c", -- 117d0
		x"00000002", -- 117d4
		x"00084a28", -- 117d8
		x"00116700", -- 117dc
		x"008c3f3c", -- 117e0
		x"00022f0e", -- 117e4
		x"4ebafbf0", -- 117e8
		x"6000007e", -- 117ec
		x"3f3cfffc", -- 117f0
		x"2f0e4eba", -- 117f4
		x"fc986000", -- 117f8
		x"0070206e", -- 117fc
		x"ffe24aa8", -- 11800
		x"00226f2e", -- 11804
		x"20280022", -- 11808
		x"e7802170", -- 1180c
		x"081e0004", -- 11810
		x"2d700822", -- 11814
		x"fffa53a8", -- 11818
		x"00224a28", -- 1181c
		x"0011670a", -- 11820
		x"3f3c0002", -- 11824
		x"2f0e4eba", -- 11828
		x"fbae2f0e", -- 1182c
		x"4ebafcbc", -- 11830
		x"6036206e", -- 11834
		x"ffde3f28", -- 11838
		x"00026026", -- 1183c
		x"422effff", -- 11840
		x"206effde", -- 11844
		x"226effe2", -- 11848
		x"30280002", -- 1184c
		x"48c02340", -- 11850
		x"00086014", -- 11854
		x"206effde", -- 11858
		x"3f280002", -- 1185c
		x"60043f3c", -- 11860
		x"ffff2f0e", -- 11864
		x"4ebafc26", -- 11868
		x"4a2effff", -- 1186c
		x"6600fd9a", -- 11870
		x"4e5e2e9f", -- 11874
		x"4e754e75", -- 11878
		x"4e750000", -- 1187c
		x"4e56fffc", -- 11880
		x"2d6e000a", -- 11884
		x"fffc206e", -- 11888
		x"fffc4a68", -- 1188c
		x"00306600", -- 11890
		x"0008316e", -- 11894
		x"00080030", -- 11898
		x"4e5e205f", -- 1189c
		x"5c4f4ed0", -- 118a0
		x"4e750000", -- 118a4
		x"4e560000", -- 118a8
		x"23fc0000", -- 118ac
		x"00010088", -- 118b0
		x"00044e5e", -- 118b4
		x"4e750000", -- 118b8
		x"4e560000", -- 118bc
		x"42b90088", -- 118c0
		x"00044e5e", -- 118c4
		x"4e750000", -- 118c8
		x"4e560000", -- 118cc
		x"7001b0b9", -- 118d0
		x"00880004", -- 118d4
		x"66000020", -- 118d8
		x"52b90088", -- 118dc
		x"00082039", -- 118e0
		x"00880008", -- 118e4
		x"e58041f9", -- 118e8
		x"00880004", -- 118ec
		x"d0fc0004", -- 118f0
		x"21ae0008", -- 118f4
		x"08004e5e", -- 118f8
		x"2e9f4e75", -- 118fc
		x"00004e56", -- 11900
		x"fff22079", -- 11904
		x"fffffed4", -- 11908
		x"2d680010", -- 1190c
		x"fffa206e", -- 11910
		x"fffa41e8", -- 11914
		x"00162d48", -- 11918
		x"fff6206e", -- 1191c
		x"fff6317c", -- 11920
		x"ffff0004", -- 11924
		x"42104228", -- 11928
		x"00014228", -- 1192c
		x"0002316e", -- 11930
		x"00080006", -- 11934
		x"2f3c0001", -- 11938
		x"0000302e", -- 1193c
		x"000848c0", -- 11940
		x"2f004eb9", -- 11944
		x"000081b0", -- 11948
		x"06970060", -- 1194c
		x"0000206e", -- 11950
		x"fff6215f", -- 11954
		x"00082268", -- 11958
		x"00081029", -- 1195c
		x"00010200", -- 11960
		x"001f7200", -- 11964
		x"12003141", -- 11968
		x"000c43e8", -- 1196c
		x"000e2d49", -- 11970
		x"fff23d7c", -- 11974
		x"fffffffe", -- 11978
		x"526efffe", -- 1197c
		x"206efff2", -- 11980
		x"302efffe", -- 11984
		x"48c0e580", -- 11988
		x"42b00800", -- 1198c
		x"302efffe", -- 11990
		x"48c0e580", -- 11994
		x"31bc0001", -- 11998
		x"0820302e", -- 1199c
		x"fffe48c0", -- 119a0
		x"e58011bc", -- 119a4
		x"ff000823", -- 119a8
		x"0c6e0007", -- 119ac
		x"fffe6dc8", -- 119b0
		x"206efff6", -- 119b4
		x"226efff2", -- 119b8
		x"23680008", -- 119bc
		x"00402368", -- 119c0
		x"00080044", -- 119c4
		x"06a90000", -- 119c8
		x"00200044", -- 119cc
		x"24690040", -- 119d0
		x"102a0003", -- 119d4
		x"e8880280", -- 119d8
		x"00000003", -- 119dc
		x"56803340", -- 119e0
		x"0048336e", -- 119e4
		x"0008004a", -- 119e8
		x"4229004c", -- 119ec
		x"237cffff", -- 119f0
		x"ffff004e", -- 119f4
		x"4e5e205f", -- 119f8
		x"544f4ed0", -- 119fc
		x"00004e56", -- 11a00
		x"fff842ae", -- 11a04
		x"000a2079", -- 11a08
		x"fffffed4", -- 11a0c
		x"2d680010", -- 11a10
		x"fffc206e", -- 11a14
		x"fffc41e8", -- 11a18
		x"00162d48", -- 11a1c
		x"fff8206e", -- 11a20
		x"fff8302e", -- 11a24
		x"0008b068", -- 11a28
		x"00066600", -- 11a2c
		x"00147007", -- 11a30
		x"b068000c", -- 11a34
		x"6600000a", -- 11a38
		x"43e8000e", -- 11a3c
		x"2d49000a", -- 11a40
		x"4e5e205f", -- 11a44
		x"544f4ed0", -- 11a48
		x"00004e56", -- 11a4c
		x"fff42079", -- 11a50
		x"fffffed4", -- 11a54
		x"2d680010", -- 11a58
		x"fff8206e", -- 11a5c
		x"fff841e8", -- 11a60
		x"00162d48", -- 11a64
		x"fff4206e", -- 11a68
		x"fff443e8", -- 11a6c
		x"000e2d49", -- 11a70
		x"fffc206e", -- 11a74
		x"fffc4cae", -- 11a78
		x"1e00000a", -- 11a7c
		x"48a81e00", -- 11a80
		x"00524e5e", -- 11a84
		x"205fdefc", -- 11a88
		x"000a4ed0", -- 11a8c
		x"00004e56", -- 11a90
		x"00002079", -- 11a94
		x"fffffed4", -- 11a98
		x"08280005", -- 11a9c
		x"000b56c0", -- 11aa0
		x"44004a00", -- 11aa4
		x"67000042", -- 11aa8
		x"2f2dfff6", -- 11aac
		x"2f0e487a", -- 11ab0
		x"002a2b4f", -- 11ab4
		x"fff64ab9", -- 11ab8
		x"00500010", -- 11abc
		x"57c00200", -- 11ac0
		x"00011d40", -- 11ac4
		x"00081d7c", -- 11ac8
		x"00010008", -- 11acc
		x"2b6f0008", -- 11ad0
		x"fff6defc", -- 11ad4
		x"000c4efa", -- 11ad8
		x"000c2c5f", -- 11adc
		x"2b5ffff6", -- 11ae0
		x"422e0008", -- 11ae4
		x"60000006", -- 11ae8
		x"422e0008", -- 11aec
		x"422e0008", -- 11af0
		x"4e5e4e75", -- 11af4
		x"00004e56", -- 11af8
		x"fff82079", -- 11afc
		x"fffffed4", -- 11b00
		x"08280005", -- 11b04
		x"000b56c0", -- 11b08
		x"44004a00", -- 11b0c
		x"6700005e", -- 11b10
		x"2079ffff", -- 11b14
		x"fed42d68", -- 11b18
		x"0010fffc", -- 11b1c
		x"206efffc", -- 11b20
		x"41e80016", -- 11b24
		x"2d48fff8", -- 11b28
		x"206efff8", -- 11b2c
		x"317cffff", -- 11b30
		x"00044a28", -- 11b34
		x"00016600", -- 11b38
		x"000a4268", -- 11b3c
		x"00046000", -- 11b40
		x"0014206e", -- 11b44
		x"fff84a28", -- 11b48
		x"00026600", -- 11b4c
		x"0008317c", -- 11b50
		x"00010004", -- 11b54
		x"206efff8", -- 11b58
		x"30280004", -- 11b5c
		x"11bc0001", -- 11b60
		x"00013028", -- 11b64
		x"000448c0", -- 11b68
		x"2d40000a", -- 11b6c
		x"2d7cffff", -- 11b70
		x"ffff000a", -- 11b74
		x"4e5e205f", -- 11b78
		x"544f4ed0", -- 11b7c
		x"00004e56", -- 11b80
		x"ffe0206e", -- 11b84
		x"000c4a10", -- 11b88
		x"67000050", -- 11b8c
		x"206e000c", -- 11b90
		x"4210558f", -- 11b94
		x"4ebafef8", -- 11b98
		x"4a1f6700", -- 11b9c
		x"003e206e", -- 11ba0
		x"00082d68", -- 11ba4
		x"0010ffec", -- 11ba8
		x"202effec", -- 11bac
		x"02800000", -- 11bb0
		x"00034a80", -- 11bb4
		x"66000024", -- 11bb8
		x"206e0008", -- 11bbc
		x"2d680014", -- 11bc0
		x"ffec202e", -- 11bc4
		x"ffec0280", -- 11bc8
		x"00000003", -- 11bcc
		x"4a806600", -- 11bd0
		x"000a206e", -- 11bd4
		x"000c10bc", -- 11bd8
		x"00012f2e", -- 11bdc
		x"0010206e", -- 11be0
		x"000c1f10", -- 11be4
		x"4eb90001", -- 11be8
		x"1d942d7c", -- 11bec
		x"00500000", -- 11bf0
		x"fffc206e", -- 11bf4
		x"000c4a10", -- 11bf8
		x"67000098", -- 11bfc
		x"2d6efffc", -- 11c00
		x"fff006ae", -- 11c04
		x"00000010", -- 11c08
		x"fff0202e", -- 11c0c
		x"00105280", -- 11c10
		x"e1802d6e", -- 11c14
		x"fffcfff4", -- 11c18
		x"d1aefff4", -- 11c1c
		x"2d6efff0", -- 11c20
		x"ffe82d6e", -- 11c24
		x"fff4ffe4", -- 11c28
		x"2d6e0008", -- 11c2c
		x"ffe0206e", -- 11c30
		x"ffe80228", -- 11c34
		x"fffc0005", -- 11c38
		x"70008128", -- 11c3c
		x"00050228", -- 11c40
		x"00f30005", -- 11c44
		x"7002e588", -- 11c48
		x"81280005", -- 11c4c
		x"226effe0", -- 11c50
		x"246effe4", -- 11c54
		x"24a90010", -- 11c58
		x"23690014", -- 11c5c
		x"000c2029", -- 11c60
		x"00146c02", -- 11c64
		x"5680e480", -- 11c68
		x"53802540", -- 11c6c
		x"0004266e", -- 11c70
		x"00087001", -- 11c74
		x"b0536600", -- 11c78
		x"000c357c", -- 11c7c
		x"810a0008", -- 11c80
		x"6000000c", -- 11c84
		x"206effe4", -- 11c88
		x"317c810e", -- 11c8c
		x"00086000", -- 11c90
		x"008e202e", -- 11c94
		x"0010e780", -- 11c98
		x"2d6efffc", -- 11c9c
		x"fff8d1ae", -- 11ca0
		x"fff82d6e", -- 11ca4
		x"fff8ffe8", -- 11ca8
		x"2d6e0008", -- 11cac
		x"ffe4206e", -- 11cb0
		x"ffe4226e", -- 11cb4
		x"ffe822a8", -- 11cb8
		x"00100ca8", -- 11cbc
		x"00020000", -- 11cc0
		x"00146d00", -- 11cc4
		x"0016217c", -- 11cc8
		x"00020000", -- 11ccc
		x"000c2d7c", -- 11cd0
		x"0000ffff", -- 11cd4
		x"ffec6000", -- 11cd8
		x"001c206e", -- 11cdc
		x"ffe42168", -- 11ce0
		x"0014000c", -- 11ce4
		x"20280014", -- 11ce8
		x"6c025280", -- 11cec
		x"e2805380", -- 11cf0
		x"2d40ffec", -- 11cf4
		x"206effe8", -- 11cf8
		x"316effee", -- 11cfc
		x"0004226e", -- 11d00
		x"00087001", -- 11d04
		x"b0516600", -- 11d08
		x"000c317c", -- 11d0c
		x"810a0006", -- 11d10
		x"6000000c", -- 11d14
		x"206effe8", -- 11d18
		x"317c810e", -- 11d1c
		x"00064e5e", -- 11d20
		x"205fdefc", -- 11d24
		x"000c4ed0", -- 11d28
		x"00004e56", -- 11d2c
		x"fff84a2e", -- 11d30
		x"000c6700", -- 11d34
		x"0014202e", -- 11d38
		x"000e5280", -- 11d3c
		x"e1805080", -- 11d40
		x"2d40fff8", -- 11d44
		x"6000000e", -- 11d48
		x"202e000e", -- 11d4c
		x"e7805c80", -- 11d50
		x"2d40fff8", -- 11d54
		x"2d7c0050", -- 11d58
		x"0000fffc", -- 11d5c
		x"202efff8", -- 11d60
		x"d1aefffc", -- 11d64
		x"206e0008", -- 11d68
		x"7001b050", -- 11d6c
		x"6600000e", -- 11d70
		x"206efffc", -- 11d74
		x"30bc810a", -- 11d78
		x"6000000a", -- 11d7c
		x"206efffc", -- 11d80
		x"30bc810e", -- 11d84
		x"4e5e205f", -- 11d88
		x"defc000a", -- 11d8c
		x"4ed00000", -- 11d90
		x"4e56fffa", -- 11d94
		x"4a2e0008", -- 11d98
		x"67000036", -- 11d9c
		x"2d7c0050", -- 11da0
		x"0000fffa", -- 11da4
		x"06ae0000", -- 11da8
		x"0010fffa", -- 11dac
		x"4aae000a", -- 11db0
		x"66000010", -- 11db4
		x"206efffa", -- 11db8
		x"08e80004", -- 11dbc
		x"00056000", -- 11dc0
		x"000c206e", -- 11dc4
		x"fffa08e8", -- 11dc8
		x"00050005", -- 11dcc
		x"60000018", -- 11dd0
		x"202e000a", -- 11dd4
		x"e78041f9", -- 11dd8
		x"00500000", -- 11ddc
		x"48700800", -- 11de0
		x"205f3d50", -- 11de4
		x"fffe4e5e", -- 11de8
		x"205f5c4f", -- 11dec
		x"4ed00000", -- 11df0
		x"4e56ffe8", -- 11df4
		x"1d7c0001", -- 11df8
		x"00122d7c", -- 11dfc
		x"00500000", -- 11e00
		x"fffc4a2e", -- 11e04
		x"000c6700", -- 11e08
		x"0080202e", -- 11e0c
		x"000e5280", -- 11e10
		x"e1802d6e", -- 11e14
		x"fffcfff8", -- 11e18
		x"d1aefff8", -- 11e1c
		x"2d6efff8", -- 11e20
		x"ffe8202e", -- 11e24
		x"00086c02", -- 11e28
		x"5680e480", -- 11e2c
		x"53802d40", -- 11e30
		x"fff4206e", -- 11e34
		x"ffe82028", -- 11e38
		x"0004b0ae", -- 11e3c
		x"fff46700", -- 11e40
		x"00442f3c", -- 11e44
		x"000f4240", -- 11e48
		x"4eb90001", -- 11e4c
		x"4b16206e", -- 11e50
		x"ffe82028", -- 11e54
		x"0004b0ae", -- 11e58
		x"fff457c0", -- 11e5c
		x"67000012", -- 11e60
		x"558f4eb9", -- 11e64
		x"00014b30", -- 11e68
		x"101f6600", -- 11e6c
		x"000460de", -- 11e70
		x"206effe8", -- 11e74
		x"20280004", -- 11e78
		x"b0aefff4", -- 11e7c
		x"67000006", -- 11e80
		x"422e0012", -- 11e84
		x"60000086", -- 11e88
		x"202e000e", -- 11e8c
		x"e7802d6e", -- 11e90
		x"fffcfff0", -- 11e94
		x"d1aefff0", -- 11e98
		x"2d6efff0", -- 11e9c
		x"ffe8202e", -- 11ea0
		x"00086c02", -- 11ea4
		x"5280e280", -- 11ea8
		x"53800280", -- 11eac
		x"0000ffff", -- 11eb0
		x"2d40ffec", -- 11eb4
		x"206effe8", -- 11eb8
		x"70003028", -- 11ebc
		x"0004b0ae", -- 11ec0
		x"ffec6700", -- 11ec4
		x"00482f3c", -- 11ec8
		x"000f4240", -- 11ecc
		x"4eb90001", -- 11ed0
		x"4b16206e", -- 11ed4
		x"ffe87000", -- 11ed8
		x"30280004", -- 11edc
		x"b0aeffec", -- 11ee0
		x"57c06700", -- 11ee4
		x"0012558f", -- 11ee8
		x"4eb90001", -- 11eec
		x"4b30101f", -- 11ef0
		x"66000004", -- 11ef4
		x"60dc206e", -- 11ef8
		x"ffe87000", -- 11efc
		x"30280004", -- 11f00
		x"b0aeffec", -- 11f04
		x"67000006", -- 11f08
		x"422e0012", -- 11f0c
		x"2f2e000e", -- 11f10
		x"1f2e000c", -- 11f14
		x"4ebafe7a", -- 11f18
		x"4e5e205f", -- 11f1c
		x"defc000a", -- 11f20
		x"4ed00000", -- 11f24
		x"4e56fff8", -- 11f28
		x"2079ffff", -- 11f2c
		x"fed42d68", -- 11f30
		x"0010fffc", -- 11f34
		x"206efffc", -- 11f38
		x"41e80016", -- 11f3c
		x"2d48fff8", -- 11f40
		x"206efff8", -- 11f44
		x"30280004", -- 11f48
		x"42300001", -- 11f4c
		x"4e5e205f", -- 11f50
		x"544f4ed0", -- 11f54
		x"4e750000", -- 11f58
		x"00080000", -- 11f5c
		x"00080000", -- 11f60
		x"00070000", -- 11f64
		x"00090000", -- 11f68
		x"00030000", -- 11f6c
		x"00010000", -- 11f70
		x"00060000", -- 11f74
		x"00050000", -- 11f78
		x"4e56fff6", -- 11f7c
		x"2d6e000c", -- 11f80
		x"fffa206e", -- 11f84
		x"fffa2268", -- 11f88
		x"00482d69", -- 11f8c
		x"0044fff6", -- 11f90
		x"206efff6", -- 11f94
		x"1d68000b", -- 11f98
		x"ffff1028", -- 11f9c
		x"000de888", -- 11fa0
		x"02800000", -- 11fa4
		x"000f6600", -- 11fa8
		x"002e082e", -- 11fac
		x"0003ffff", -- 11fb0
		x"56c04400", -- 11fb4
		x"4a006700", -- 11fb8
		x"0010226e", -- 11fbc
		x"000822bc", -- 11fc0
		x"00000004", -- 11fc4
		x"6000000c", -- 11fc8
		x"206e0008", -- 11fcc
		x"20bc0000", -- 11fd0
		x"00036000", -- 11fd4
		x"0048206e", -- 11fd8
		x"fffa7001", -- 11fdc
		x"b068002c", -- 11fe0
		x"67000010", -- 11fe4
		x"226e0008", -- 11fe8
		x"22bc0000", -- 11fec
		x"00046000", -- 11ff0
		x"002c102e", -- 11ff4
		x"ffff0280", -- 11ff8
		x"00000007", -- 11ffc
		x"e580206e", -- 12000
		x"000843fa", -- 12004
		x"ff5220b1", -- 12008
		x"0800206e", -- 1200c
		x"00087001", -- 12010
		x"b0906600", -- 12014
		x"00081d7c", -- 12018
		x"00ffffff", -- 1201c
		x"206efff6", -- 12020
		x"102effff", -- 12024
		x"b028000b", -- 12028
		x"6600ff66", -- 1202c
		x"4e5e205f", -- 12030
		x"504f4ed0", -- 12034
		x"00004e56", -- 12038
		x"0000206e", -- 1203c
		x"000c3f10", -- 12040
		x"4eb90001", -- 12044
		x"227e206e", -- 12048
		x"00084290", -- 1204c
		x"4e5e205f", -- 12050
		x"504f4ed0", -- 12054
		x"00004e56", -- 12058
		x"0000206e", -- 1205c
		x"000c3f10", -- 12060
		x"4eb90001", -- 12064
		x"236a206e", -- 12068
		x"00084290", -- 1206c
		x"4e5e205f", -- 12070
		x"504f4ed0", -- 12074
		x"00004e56", -- 12078
		x"ffee206e", -- 1207c
		x"000c2068", -- 12080
		x"00482d68", -- 12084
		x"0044fff6", -- 12088
		x"206efff6", -- 1208c
		x"598f7000", -- 12090
		x"1028001b", -- 12094
		x"2f002f3c", -- 12098
		x"00000008", -- 1209c
		x"2d48fff2", -- 120a0
		x"4eb90001", -- 120a4
		x"4b5a206e", -- 120a8
		x"fff2598f", -- 120ac
		x"70001028", -- 120b0
		x"00192f00", -- 120b4
		x"2f3c0000", -- 120b8
		x"00102d48", -- 120bc
		x"ffee4eb9", -- 120c0
		x"00014b5a", -- 120c4
		x"206effee", -- 120c8
		x"201fd09f", -- 120cc
		x"72001228", -- 120d0
		x"001dd081", -- 120d4
		x"d0bc0000", -- 120d8
		x"04002d40", -- 120dc
		x"fffc0228", -- 120e0
		x"ff1f0005", -- 120e4
		x"7003eb88", -- 120e8
		x"81280005", -- 120ec
		x"206efff6", -- 120f0
		x"1028000b", -- 120f4
		x"02800000", -- 120f8
		x"00077206", -- 120fc
		x"b2806700", -- 12100
		x"01344aae", -- 12104
		x"fffc6f00", -- 12108
		x"012c2f3c", -- 1210c
		x"000f4240", -- 12110
		x"4eb90001", -- 12114
		x"4b16206e", -- 12118
		x"fff60828", -- 1211c
		x"0007000b", -- 12120
		x"56c04400", -- 12124
		x"66000012", -- 12128
		x"558f4eb9", -- 1212c
		x"00014b30", -- 12130
		x"101f6600", -- 12134
		x"000460de", -- 12138
		x"206efff6", -- 1213c
		x"08280007", -- 12140
		x"000b56c0", -- 12144
		x"44000840", -- 12148
		x"00006700", -- 1214c
		x"001a1028", -- 12150
		x"000b0280", -- 12154
		x"00000007", -- 12158
		x"7206b280", -- 1215c
		x"57c06700", -- 12160
		x"00066000", -- 12164
		x"00066000", -- 12168
		x"00cc206e", -- 1216c
		x"fff61028", -- 12170
		x"000b0228", -- 12174
		x"00f80011", -- 12178
		x"02000007", -- 1217c
		x"81280011", -- 12180
		x"08280000", -- 12184
		x"000b56c0", -- 12188
		x"44004a00", -- 1218c
		x"6700004a", -- 12190
		x"0228001f", -- 12194
		x"00057007", -- 12198
		x"eb888128", -- 1219c
		x"0005206e", -- 121a0
		x"fff60828", -- 121a4
		x"0007000b", -- 121a8
		x"56c04400", -- 121ac
		x"08400000", -- 121b0
		x"67000018", -- 121b4
		x"1028000b", -- 121b8
		x"02800000", -- 121bc
		x"00077206", -- 121c0
		x"b28057c0", -- 121c4
		x"67000004", -- 121c8
		x"60d4206e", -- 121cc
		x"fff61d68", -- 121d0
		x"0017fffb", -- 121d4
		x"60000044", -- 121d8
		x"206efff6", -- 121dc
		x"42280017", -- 121e0
		x"0228001f", -- 121e4
		x"00057007", -- 121e8
		x"eb888128", -- 121ec
		x"0005206e", -- 121f0
		x"fff60828", -- 121f4
		x"0007000b", -- 121f8
		x"56c04400", -- 121fc
		x"08400000", -- 12200
		x"67000018", -- 12204
		x"1028000b", -- 12208
		x"02800000", -- 1220c
		x"00077206", -- 12210
		x"b28057c0", -- 12214
		x"67000004", -- 12218
		x"60d4206e", -- 1221c
		x"fff60228", -- 12220
		x"ff1f0005", -- 12224
		x"7006eb88", -- 12228
		x"81280005", -- 1222c
		x"53aefffc", -- 12230
		x"6000feba", -- 12234
		x"206efff6", -- 12238
		x"1028000b", -- 1223c
		x"02800000", -- 12240
		x"00077206", -- 12244
		x"b2806700", -- 12248
		x"001e226e", -- 1224c
		x"000822bc", -- 12250
		x"00000001", -- 12254
		x"2f2e000c", -- 12258
		x"3f3c000b", -- 1225c
		x"4eb90001", -- 12260
		x"18806000", -- 12264
		x"000c206e", -- 12268
		x"000820bc", -- 1226c
		x"00000006", -- 12270
		x"4e5e205f", -- 12274
		x"504f4ed0", -- 12278
		x"00004e56", -- 1227c
		x"fff0598f", -- 12280
		x"3f2e0008", -- 12284
		x"4eb90001", -- 12288
		x"1a022d5f", -- 1228c
		x"fffc2d6e", -- 12290
		x"fffcfff8", -- 12294
		x"206efff8", -- 12298
		x"2d680044", -- 1229c
		x"fff42d68", -- 122a0
		x"0040fff0", -- 122a4
		x"226efff0", -- 122a8
		x"137cff00", -- 122ac
		x"000108a9", -- 122b0
		x"00070003", -- 122b4
		x"246efff4", -- 122b8
		x"157cff00", -- 122bc
		x"0003157c", -- 122c0
		x"ffc00003", -- 122c4
		x"2f3c0000", -- 122c8
		x"03e84eb9", -- 122cc
		x"00014b10", -- 122d0
		x"206efff0", -- 122d4
		x"10280007", -- 122d8
		x"02800000", -- 122dc
		x"00077207", -- 122e0
		x"9280226e", -- 122e4
		x"fff41341", -- 122e8
		x"0001137c", -- 122ec
		x"00000005", -- 122f0
		x"137c0000", -- 122f4
		x"0007137c", -- 122f8
		x"00000011", -- 122fc
		x"42290017", -- 12300
		x"42290019", -- 12304
		x"4229001b", -- 12308
		x"4229001d", -- 1230c
		x"137c0000", -- 12310
		x"000b1369", -- 12314
		x"00090009", -- 12318
		x"08280003", -- 1231c
		x"000756c0", -- 12320
		x"44004a00", -- 12324
		x"6700000c", -- 12328
		x"137c0099", -- 1232c
		x"00036000", -- 12330
		x"000c206e", -- 12334
		x"fff4117c", -- 12338
		x"ff910003", -- 1233c
		x"206efff4", -- 12340
		x"08a80007", -- 12344
		x"0003226e", -- 12348
		x"fff0137c", -- 1234c
		x"ff010007", -- 12350
		x"2f3c0000", -- 12354
		x"03e84eb9", -- 12358
		x"00014b10", -- 1235c
		x"4e5e205f", -- 12360
		x"544f4ed0", -- 12364
		x"00004e56", -- 12368
		x"ffec598f", -- 1236c
		x"3f2e0008", -- 12370
		x"4eb90001", -- 12374
		x"1a022d5f", -- 12378
		x"fffc2d6e", -- 1237c
		x"fffcfff4", -- 12380
		x"206efff4", -- 12384
		x"2d680040", -- 12388
		x"fff02d68", -- 1238c
		x"0044ffec", -- 12390
		x"226efff0", -- 12394
		x"08a90007", -- 12398
		x"0003246e", -- 1239c
		x"ffec157c", -- 123a0
		x"ff000003", -- 123a4
		x"157cff10", -- 123a8
		x"00052f3c", -- 123ac
		x"000003e8", -- 123b0
		x"4eb90001", -- 123b4
		x"4b10206e", -- 123b8
		x"ffec117c", -- 123bc
		x"ffc00003", -- 123c0
		x"2f3c0000", -- 123c4
		x"03e84eb9", -- 123c8
		x"00014b10", -- 123cc
		x"206effec", -- 123d0
		x"08a80007", -- 123d4
		x"0003226e", -- 123d8
		x"fff0137c", -- 123dc
		x"ff010007", -- 123e0
		x"2d7cffff", -- 123e4
		x"fffffff8", -- 123e8
		x"52aefff8", -- 123ec
		x"206efff4", -- 123f0
		x"202efff8", -- 123f4
		x"e58031bc", -- 123f8
		x"00010820", -- 123fc
		x"0cae0000", -- 12400
		x"0007fff8", -- 12404
		x"6de22f3c", -- 12408
		x"001e8480", -- 1240c
		x"4eb90001", -- 12410
		x"4b104e5e", -- 12414
		x"205f544f", -- 12418
		x"4ed00000", -- 1241c
		x"4e560000", -- 12420
		x"206e0008", -- 12424
		x"20680048", -- 12428
		x"2d680040", -- 1242c
		x"000c4e5e", -- 12430
		x"2e9f4e75", -- 12434
		x"00004e56", -- 12438
		x"0000206e", -- 1243c
		x"00082068", -- 12440
		x"00482d68", -- 12444
		x"0044000c", -- 12448
		x"4e5e2e9f", -- 1244c
		x"4e750000", -- 12450
		x"4e56fff8", -- 12454
		x"206e0012", -- 12458
		x"20680048", -- 1245c
		x"2d680044", -- 12460
		x"fff8206e", -- 12464
		x"fff81168", -- 12468
		x"00090009", -- 1246c
		x"117c0000", -- 12470
		x"00074a2e", -- 12474
		x"000a6700", -- 12478
		x"00227006", -- 1247c
		x"b06e000c", -- 12480
		x"66000018", -- 12484
		x"206efff8", -- 12488
		x"0228ff1f", -- 1248c
		x"00057003", -- 12490
		x"eb888128", -- 12494
		x"00056000", -- 12498
		x"0014206e", -- 1249c
		x"fff80228", -- 124a0
		x"ff1f0005", -- 124a4
		x"7002eb88", -- 124a8
		x"81280005", -- 124ac
		x"206efff8", -- 124b0
		x"08280007", -- 124b4
		x"000b56c0", -- 124b8
		x"44004a00", -- 124bc
		x"6600005e", -- 124c0
		x"1028000b", -- 124c4
		x"02800000", -- 124c8
		x"0007322e", -- 124cc
		x"000c48c1", -- 124d0
		x"b0816600", -- 124d4
		x"00482f3c", -- 124d8
		x"000f4240", -- 124dc
		x"4eb90001", -- 124e0
		x"4b16206e", -- 124e4
		x"fff80828", -- 124e8
		x"0007000b", -- 124ec
		x"56c04400", -- 124f0
		x"6600002a", -- 124f4
		x"1028000b", -- 124f8
		x"02800000", -- 124fc
		x"0007322e", -- 12500
		x"000c48c1", -- 12504
		x"b08156c0", -- 12508
		x"66000012", -- 1250c
		x"558f4eb9", -- 12510
		x"00014b30", -- 12514
		x"101f6600", -- 12518
		x"000460c6", -- 1251c
		x"206efff8", -- 12520
		x"08280007", -- 12524
		x"000b56c0", -- 12528
		x"44000840", -- 1252c
		x"00006700", -- 12530
		x"001e1028", -- 12534
		x"000b0280", -- 12538
		x"00000007", -- 1253c
		x"322e000c", -- 12540
		x"48c1b081", -- 12544
		x"56c06600", -- 12548
		x"00066000", -- 1254c
		x"000a422e", -- 12550
		x"00166000", -- 12554
		x"00f6206e", -- 12558
		x"fff80228", -- 1255c
		x"fff80011", -- 12560
		x"302e000c", -- 12564
		x"81280011", -- 12568
		x"08280000", -- 1256c
		x"000b56c0", -- 12570
		x"44004a00", -- 12574
		x"67000046", -- 12578
		x"0228001f", -- 1257c
		x"00057007", -- 12580
		x"eb888128", -- 12584
		x"0005206e", -- 12588
		x"fff80828", -- 1258c
		x"0007000b", -- 12590
		x"56c04400", -- 12594
		x"08400000", -- 12598
		x"6700000e", -- 1259c
		x"4a280009", -- 125a0
		x"56c06600", -- 125a4
		x"000460de", -- 125a8
		x"206efff8", -- 125ac
		x"226e000e", -- 125b0
		x"70001028", -- 125b4
		x"00173280", -- 125b8
		x"60000040", -- 125bc
		x"206e000e", -- 125c0
		x"226efff8", -- 125c4
		x"13680001", -- 125c8
		x"00170229", -- 125cc
		x"001f0005", -- 125d0
		x"7007eb88", -- 125d4
		x"81290005", -- 125d8
		x"206efff8", -- 125dc
		x"08280007", -- 125e0
		x"000b56c0", -- 125e4
		x"44000840", -- 125e8
		x"00006700", -- 125ec
		x"000e4a28", -- 125f0
		x"000956c0", -- 125f4
		x"66000004", -- 125f8
		x"60de206e", -- 125fc
		x"fff84a28", -- 12600
		x"00096600", -- 12604
		x"00301d7c", -- 12608
		x"00010016", -- 1260c
		x"7007b06e", -- 12610
		x"000c6600", -- 12614
		x"001c4a2e", -- 12618
		x"00086700", -- 1261c
		x"0014206e", -- 12620
		x"fff80228", -- 12624
		x"ff1f0005", -- 12628
		x"7003eb88", -- 1262c
		x"81280005", -- 12630
		x"60000006", -- 12634
		x"422e0016", -- 12638
		x"206efff8", -- 1263c
		x"0228ff1f", -- 12640
		x"00057006", -- 12644
		x"eb888128", -- 12648
		x"00054a2e", -- 1264c
		x"000a6600", -- 12650
		x"008c206e", -- 12654
		x"fff84a28", -- 12658
		x"00096600", -- 1265c
		x"0080206e", -- 12660
		x"fff81028", -- 12664
		x"000b0280", -- 12668
		x"00000007", -- 1266c
		x"322e000c", -- 12670
		x"48c1b280", -- 12674
		x"66000066", -- 12678
		x"2f3c000f", -- 1267c
		x"42404eb9", -- 12680
		x"00014b16", -- 12684
		x"206efff8", -- 12688
		x"1028000b", -- 1268c
		x"02800000", -- 12690
		x"0007322e", -- 12694
		x"000c48c1", -- 12698
		x"b28056c0", -- 1269c
		x"66000012", -- 126a0
		x"558f4eb9", -- 126a4
		x"00014b30", -- 126a8
		x"101f6600", -- 126ac
		x"000460d4", -- 126b0
		x"206efff8", -- 126b4
		x"1028000b", -- 126b8
		x"02800000", -- 126bc
		x"0007322e", -- 126c0
		x"000c48c1", -- 126c4
		x"b2806600", -- 126c8
		x"0014422e", -- 126cc
		x"00162f2e", -- 126d0
		x"00123f3c", -- 126d4
		x"000b4eb9", -- 126d8
		x"00011880", -- 126dc
		x"206efff8", -- 126e0
		x"11680009", -- 126e4
		x"00094e5e", -- 126e8
		x"205fdefc", -- 126ec
		x"000e4ed0", -- 126f0
		x"00004e56", -- 126f4
		x"ffea1d7c", -- 126f8
		x"0001000c", -- 126fc
		x"206e0008", -- 12700
		x"41e80044", -- 12704
		x"2d48fff6", -- 12708
		x"206efff6", -- 1270c
		x"2d680004", -- 12710
		x"fff2226e", -- 12714
		x"fff22d69", -- 12718
		x"0040ffee", -- 1271c
		x"2d690044", -- 12720
		x"ffea246e", -- 12724
		x"ffee082a", -- 12728
		x"00050001", -- 1272c
		x"56c04400", -- 12730
		x"08400000", -- 12734
		x"02000001", -- 12738
		x"1340004d", -- 1273c
		x"08aa0000", -- 12740
		x"000308aa", -- 12744
		x"00010003", -- 12748
		x"2f29004e", -- 1274c
		x"4869004d", -- 12750
		x"48680014", -- 12754
		x"4eb90001", -- 12758
		x"1b82206e", -- 1275c
		x"ffea117c", -- 12760
		x"ff000009", -- 12764
		x"226efff6", -- 12768
		x"137cff01", -- 1276c
		x"000e337c", -- 12770
		x"001a0010", -- 12774
		x"2d690020", -- 12778
		x"fffa202e", -- 1277c
		x"fffa6c06", -- 12780
		x"d0bc0000", -- 12784
		x"00ffe080", -- 12788
		x"6c06d0bc", -- 1278c
		x"000000ff", -- 12790
		x"e0801140", -- 12794
		x"0019202e", -- 12798
		x"fffa6c06", -- 1279c
		x"d0bc0000", -- 127a0
		x"00ffe080", -- 127a4
		x"1140001b", -- 127a8
		x"116efffd", -- 127ac
		x"001d0228", -- 127b0
		x"fff80011", -- 127b4
		x"30290014", -- 127b8
		x"81280011", -- 127bc
		x"117c0080", -- 127c0
		x"00051028", -- 127c4
		x"000de888", -- 127c8
		x"02800000", -- 127cc
		x"000f720b", -- 127d0
		x"b2806700", -- 127d4
		x"007c4a28", -- 127d8
		x"00096600", -- 127dc
		x"00742f3c", -- 127e0
		x"000f4240", -- 127e4
		x"4eb90001", -- 127e8
		x"4b16206e", -- 127ec
		x"ffea1028", -- 127f0
		x"000de888", -- 127f4
		x"02800000", -- 127f8
		x"000f720b", -- 127fc
		x"b28057c0", -- 12800
		x"6700001c", -- 12804
		x"4a280009", -- 12808
		x"56c06600", -- 1280c
		x"0012558f", -- 12810
		x"4eb90001", -- 12814
		x"4b30101f", -- 12818
		x"66000004", -- 1281c
		x"60cc206e", -- 12820
		x"ffea1028", -- 12824
		x"000de888", -- 12828
		x"02800000", -- 1282c
		x"000f720b", -- 12830
		x"b2806700", -- 12834
		x"001c4a28", -- 12838
		x"00096600", -- 1283c
		x"0014422e", -- 12840
		x"000c2f2e", -- 12844
		x"00083f3c", -- 12848
		x"000c4eb9", -- 1284c
		x"00011880", -- 12850
		x"206effea", -- 12854
		x"1028000d", -- 12858
		x"e8880280", -- 1285c
		x"0000000f", -- 12860
		x"720bb280", -- 12864
		x"66000070", -- 12868
		x"4a280009", -- 1286c
		x"66000068", -- 12870
		x"1d7c0000", -- 12874
		x"ffff08ae", -- 12878
		x"0007ffff", -- 1287c
		x"206efff2", -- 12880
		x"08ae0003", -- 12884
		x"ffff1028", -- 12888
		x"004de788", -- 1288c
		x"812effff", -- 12890
		x"226efff6", -- 12894
		x"7001b069", -- 12898
		x"00146600", -- 1289c
		x"000c08ee", -- 128a0
		x"0002ffff", -- 128a4
		x"60000008", -- 128a8
		x"08ae0002", -- 128ac
		x"ffff206e", -- 128b0
		x"fff27001", -- 128b4
		x"b0a8004e", -- 128b8
		x"6600000c", -- 128bc
		x"08ee0001", -- 128c0
		x"ffff6000", -- 128c4
		x"000808ee", -- 128c8
		x"0000ffff", -- 128cc
		x"206effee", -- 128d0
		x"116effff", -- 128d4
		x"00034e5e", -- 128d8
		x"2e9f4e75", -- 128dc
		x"00004e56", -- 128e0
		x"ffe2206e", -- 128e4
		x"000c41e8", -- 128e8
		x"00442d48", -- 128ec
		x"fff2206e", -- 128f0
		x"fff243e8", -- 128f4
		x"00142d49", -- 128f8
		x"ffee2d68", -- 128fc
		x"0004ffea", -- 12900
		x"226effea", -- 12904
		x"2d690044", -- 12908
		x"ffe62d69", -- 1290c
		x"0040ffe2", -- 12910
		x"246effe2", -- 12914
		x"08aa0007", -- 12918
		x"00034228", -- 1291c
		x"000e266e", -- 12920
		x"00084293", -- 12924
		x"1d7c0001", -- 12928
		x"0010266e", -- 1292c
		x"ffe61d6b", -- 12930
		x"0009ffff", -- 12934
		x"176b0009", -- 12938
		x"00094a2b", -- 1293c
		x"000f6700", -- 12940
		x"000808ee", -- 12944
		x"0001ffff", -- 12948
		x"206effe6", -- 1294c
		x"70001028", -- 12950
		x"001be180", -- 12954
		x"72001228", -- 12958
		x"0019e181", -- 1295c
		x"e181d280", -- 12960
		x"70001028", -- 12964
		x"001dd280", -- 12968
		x"2d41fffa", -- 1296c
		x"226effee", -- 12970
		x"2029000c", -- 12974
		x"90aefffa", -- 12978
		x"2d40fff6", -- 1297c
		x"202efff6", -- 12980
		x"91a90014", -- 12984
		x"20290008", -- 12988
		x"90a90014", -- 1298c
		x"23690004", -- 12990
		x"0010d1a9", -- 12994
		x"0010082e", -- 12998
		x"0001ffff", -- 1299c
		x"56c04400", -- 129a0
		x"4a006700", -- 129a4
		x"003a08ae", -- 129a8
		x"0001ffff", -- 129ac
		x"246effea", -- 129b0
		x"2f2a004e", -- 129b4
		x"1f2a004d", -- 129b8
		x"4eb90001", -- 129bc
		x"1d94206e", -- 129c0
		x"ffe608e8", -- 129c4
		x"00060003", -- 129c8
		x"08a80006", -- 129cc
		x"00032f2e", -- 129d0
		x"000c2f2e", -- 129d4
		x"00084eba", -- 129d8
		x"f69e6000", -- 129dc
		x"005a206e", -- 129e0
		x"ffee7001", -- 129e4
		x"b0506600", -- 129e8
		x"003c558f", -- 129ec
		x"226effea", -- 129f0
		x"2f29004e", -- 129f4
		x"1f29004d", -- 129f8
		x"2f2efffa", -- 129fc
		x"4eb90001", -- 12a00
		x"1df44a1f", -- 12a04
		x"6600001a", -- 12a08
		x"2f2e000c", -- 12a0c
		x"3f3c0008", -- 12a10
		x"4eb90001", -- 12a14
		x"1880206e", -- 12a18
		x"000820bc", -- 12a1c
		x"00000001", -- 12a20
		x"60000014", -- 12a24
		x"206effea", -- 12a28
		x"2f28004e", -- 12a2c
		x"1f28004d", -- 12a30
		x"4eb90001", -- 12a34
		x"1d94082e", -- 12a38
		x"0003ffff", -- 12a3c
		x"56c04400", -- 12a40
		x"4a006700", -- 12a44
		x"001808ae", -- 12a48
		x"0003ffff", -- 12a4c
		x"206effe6", -- 12a50
		x"08e80006", -- 12a54
		x"000308a8", -- 12a58
		x"00060003", -- 12a5c
		x"082e0004", -- 12a60
		x"ffff56c0", -- 12a64
		x"44004a00", -- 12a68
		x"67000024", -- 12a6c
		x"08ae0004", -- 12a70
		x"ffff206e", -- 12a74
		x"00087001", -- 12a78
		x"b0906700", -- 12a7c
		x"0012206e", -- 12a80
		x"ffee4aa8", -- 12a84
		x"00146f00", -- 12a88
		x"0006422e", -- 12a8c
		x"00104a2e", -- 12a90
		x"ffff6700", -- 12a94
		x"002a2f2e", -- 12a98
		x"000c3f3c", -- 12a9c
		x"00044eb9", -- 12aa0
		x"00011880", -- 12aa4
		x"206e0008", -- 12aa8
		x"20bc0000", -- 12aac
		x"0001206e", -- 12ab0
		x"ffe608e8", -- 12ab4
		x"00060003", -- 12ab8
		x"08a80006", -- 12abc
		x"0003206e", -- 12ac0
		x"ffe2117c", -- 12ac4
		x"ff010007", -- 12ac8
		x"08a80001", -- 12acc
		x"000308a8", -- 12ad0
		x"00000003", -- 12ad4
		x"4e5e205f", -- 12ad8
		x"504f4ed0", -- 12adc
		x"4e754e56", -- 12ae0
		x"ffde426e", -- 12ae4
		x"fff8422e", -- 12ae8
		x"000c206e", -- 12aec
		x"000841e8", -- 12af0
		x"00442d48", -- 12af4
		x"ffee43e8", -- 12af8
		x"00142d49", -- 12afc
		x"ffea2d68", -- 12b00
		x"0004ffe6", -- 12b04
		x"226effe6", -- 12b08
		x"2d690044", -- 12b0c
		x"ffe22d69", -- 12b10
		x"0040ffde", -- 12b14
		x"246effea", -- 12b18
		x"202a0014", -- 12b1c
		x"6c06d0bc", -- 12b20
		x"000000ff", -- 12b24
		x"e0806c06", -- 12b28
		x"d0bc0000", -- 12b2c
		x"00ffe080", -- 12b30
		x"266effe2", -- 12b34
		x"17400019", -- 12b38
		x"202a0014", -- 12b3c
		x"6c06d0bc", -- 12b40
		x"000000ff", -- 12b44
		x"e0801740", -- 12b48
		x"001b176a", -- 12b4c
		x"0017001d", -- 12b50
		x"022b00f8", -- 12b54
		x"00113012", -- 12b58
		x"812b0011", -- 12b5c
		x"176b0009", -- 12b60
		x"0009177c", -- 12b64
		x"00840005", -- 12b68
		x"102b000d", -- 12b6c
		x"e8880280", -- 12b70
		x"0000000f", -- 12b74
		x"720bb280", -- 12b78
		x"67622f3c", -- 12b7c
		x"000f4240", -- 12b80
		x"4eb90001", -- 12b84
		x"4b16206e", -- 12b88
		x"ffe21028", -- 12b8c
		x"000de888", -- 12b90
		x"02800000", -- 12b94
		x"000f720b", -- 12b98
		x"b28057c0", -- 12b9c
		x"67164a28", -- 12ba0
		x"00096600", -- 12ba4
		x"01e8558f", -- 12ba8
		x"4eb90001", -- 12bac
		x"4b30101f", -- 12bb0
		x"660260d2", -- 12bb4
		x"206effe2", -- 12bb8
		x"1028000d", -- 12bbc
		x"e8880280", -- 12bc0
		x"0000000f", -- 12bc4
		x"720bb280", -- 12bc8
		x"67122f2e", -- 12bcc
		x"00083f3c", -- 12bd0
		x"00084eb9", -- 12bd4
		x"00011880", -- 12bd8
		x"60000294", -- 12bdc
		x"206effea", -- 12be0
		x"7001b050", -- 12be4
		x"6600011c", -- 12be8
		x"226effee", -- 12bec
		x"4a69003a", -- 12bf0
		x"6644226e", -- 12bf4
		x"ffe247e9", -- 12bf8
		x"000949e9", -- 12bfc
		x"000d7200", -- 12c00
		x"43e90015", -- 12c04
		x"206effea", -- 12c08
		x"24680010", -- 12c0c
		x"20280014", -- 12c10
		x"6d18600a", -- 12c14
		x"4a136612", -- 12c18
		x"031466f8", -- 12c1c
		x"14d151c8", -- 12c20
		x"fff84240", -- 12c24
		x"53806ef0", -- 12c28
		x"42802140", -- 12c2c
		x"0014214a", -- 12c30
		x"00106000", -- 12c34
		x"00cc526e", -- 12c38
		x"fff8206e", -- 12c3c
		x"ffee302e", -- 12c40
		x"fff848c0", -- 12c44
		x"d0803030", -- 12c48
		x"083848c0", -- 12c4c
		x"2d40fff4", -- 12c50
		x"670000ae", -- 12c54
		x"6d00005a", -- 12c58
		x"206effe2", -- 12c5c
		x"47e80009", -- 12c60
		x"49e8000d", -- 12c64
		x"41e80015", -- 12c68
		x"226effea", -- 12c6c
		x"24690010", -- 12c70
		x"4280242e", -- 12c74
		x"fff4600a", -- 12c78
		x"4a13660c", -- 12c7c
		x"011466f8", -- 12c80
		x"14d051ca", -- 12c84
		x"fff84282", -- 12c88
		x"2d42fff4", -- 12c8c
		x"234a0010", -- 12c90
		x"206effee", -- 12c94
		x"302efff8", -- 12c98
		x"d0403030", -- 12c9c
		x"003848c0", -- 12ca0
		x"22290014", -- 12ca4
		x"9280d282", -- 12ca8
		x"23410014", -- 12cac
		x"60000048", -- 12cb0
		x"206effe2", -- 12cb4
		x"43e80009", -- 12cb8
		x"45e8000d", -- 12cbc
		x"47e80015", -- 12cc0
		x"4280222e", -- 12cc4
		x"fff44a11", -- 12cc8
		x"660a0112", -- 12ccc
		x"66f84a13", -- 12cd0
		x"528166f6", -- 12cd4
		x"2d41fff4", -- 12cd8
		x"206effee", -- 12cdc
		x"302efff8", -- 12ce0
		x"d040226e", -- 12ce4
		x"ffea3030", -- 12ce8
		x"003848c0", -- 12cec
		x"d0a90014", -- 12cf0
		x"90812340", -- 12cf4
		x"00147003", -- 12cf8
		x"b06efff8", -- 12cfc
		x"6600ff38", -- 12d00
		x"603e226e", -- 12d04
		x"ffe247e9", -- 12d08
		x"000949e9", -- 12d0c
		x"000d7201", -- 12d10
		x"206effea", -- 12d14
		x"24680010", -- 12d18
		x"20280014", -- 12d1c
		x"6d22600c", -- 12d20
		x"4a136614", -- 12d24
		x"031466f8", -- 12d28
		x"135a0015", -- 12d2c
		x"51c8fff2", -- 12d30
		x"42405380", -- 12d34
		x"6eea4280", -- 12d38
		x"21400014", -- 12d3c
		x"214a0010", -- 12d40
		x"206effe2", -- 12d44
		x"4a280009", -- 12d48
		x"66422f3c", -- 12d4c
		x"00989680", -- 12d50
		x"4eb90001", -- 12d54
		x"4b16206e", -- 12d58
		x"ffe24a28", -- 12d5c
		x"000956c0", -- 12d60
		x"660e558f", -- 12d64
		x"4eb90001", -- 12d68
		x"4b30101f", -- 12d6c
		x"660260e6", -- 12d70
		x"206effe2", -- 12d74
		x"4a280009", -- 12d78
		x"66122f2e", -- 12d7c
		x"00083f3c", -- 12d80
		x"00084eb9", -- 12d84
		x"00011880", -- 12d88
		x"600000e4", -- 12d8c
		x"206effe2", -- 12d90
		x"1d680009", -- 12d94
		x"ffff1168", -- 12d98
		x"00090009", -- 12d9c
		x"4a28000f", -- 12da0
		x"670608ee", -- 12da4
		x"0001ffff", -- 12da8
		x"082e0001", -- 12dac
		x"ffff6730", -- 12db0
		x"08ae0001", -- 12db4
		x"ffff2f2e", -- 12db8
		x"0008486e", -- 12dbc
		x"fffa4eb9", -- 12dc0
		x"0001207a", -- 12dc4
		x"7001b0ae", -- 12dc8
		x"fffa6604", -- 12dcc
		x"600000a0", -- 12dd0
		x"206effe2", -- 12dd4
		x"08e80006", -- 12dd8
		x"000308a8", -- 12ddc
		x"00060003", -- 12de0
		x"082e0003", -- 12de4
		x"ffff674c", -- 12de8
		x"08ae0003", -- 12dec
		x"ffff206e", -- 12df0
		x"ffe27000", -- 12df4
		x"1028001b", -- 12df8
		x"e1807200", -- 12dfc
		x"12280019", -- 12e00
		x"e181e181", -- 12e04
		x"d2807000", -- 12e08
		x"1028001d", -- 12e0c
		x"d280226e", -- 12e10
		x"ffea2341", -- 12e14
		x"00142029", -- 12e18
		x"000890a9", -- 12e1c
		x"00142369", -- 12e20
		x"00040010", -- 12e24
		x"d1a90010", -- 12e28
		x"08e80006", -- 12e2c
		x"000308a8", -- 12e30
		x"00060003", -- 12e34
		x"082e0004", -- 12e38
		x"ffff6706", -- 12e3c
		x"08ae0004", -- 12e40
		x"ffff4a2e", -- 12e44
		x"ffff6720", -- 12e48
		x"206effe2", -- 12e4c
		x"08e80006", -- 12e50
		x"000308a8", -- 12e54
		x"00060003", -- 12e58
		x"2f2e0008", -- 12e5c
		x"3f3c0004", -- 12e60
		x"4eb90001", -- 12e64
		x"18806006", -- 12e68
		x"1d7c0001", -- 12e6c
		x"000c4e5e", -- 12e70
		x"2e9f4e75", -- 12e74
		x"4e750000", -- 12e78
		x"4e56fff0", -- 12e7c
		x"2d6e0008", -- 12e80
		x"fff8206e", -- 12e84
		x"fff82d68", -- 12e88
		x"0048fff4", -- 12e8c
		x"4a68002c", -- 12e90
		x"66000086", -- 12e94
		x"317c0001", -- 12e98
		x"002c4868", -- 12e9c
		x"00842f2e", -- 12ea0
		x"00084879", -- 12ea4
		x"00014bd8", -- 12ea8
		x"2f3c0000", -- 12eac
		x"000a4eb9", -- 12eb0
		x"00011354", -- 12eb4
		x"206efff8", -- 12eb8
		x"4a280036", -- 12ebc
		x"67000026", -- 12ec0
		x"2f28003c", -- 12ec4
		x"2f3c0000", -- 12ec8
		x"00064eb9", -- 12ecc
		x"000081a8", -- 12ed0
		x"2d5ffffc", -- 12ed4
		x"206efff8", -- 12ed8
		x"43e80084", -- 12edc
		x"21490040", -- 12ee0
		x"6000000e", -- 12ee4
		x"42aefffc", -- 12ee8
		x"206efff8", -- 12eec
		x"42a80038", -- 12ef0
		x"206efff8", -- 12ef4
		x"48680084", -- 12ef8
		x"2f2efffc", -- 12efc
		x"2f280038", -- 12f00
		x"4eb90001", -- 12f04
		x"1320206e", -- 12f08
		x"fff84868", -- 12f0c
		x"00841f28", -- 12f10
		x"00364eb9", -- 12f14
		x"0001133a", -- 12f18
		x"206efff8", -- 12f1c
		x"48680084", -- 12f20
		x"4eb90001", -- 12f24
		x"15d0206e", -- 12f28
		x"fff843e8", -- 12f2c
		x"00842d49", -- 12f30
		x"fff0226e", -- 12f34
		x"fff04a29", -- 12f38
		x"00106700", -- 12f3c
		x"00564a69", -- 12f40
		x"000c6c00", -- 12f44
		x"004e206e", -- 12f48
		x"fff87003", -- 12f4c
		x"b068002c", -- 12f50
		x"67000040", -- 12f54
		x"206efff8", -- 12f58
		x"317c0003", -- 12f5c
		x"002c2f2e", -- 12f60
		x"00083f3c", -- 12f64
		x"00034eb9", -- 12f68
		x"00011880", -- 12f6c
		x"206efff0", -- 12f70
		x"226efff8", -- 12f74
		x"3368000c", -- 12f78
		x"004e3368", -- 12f7c
		x"000e0050", -- 12f80
		x"3f114aa9", -- 12f84
		x"007a6704", -- 12f88
		x"2f29007a", -- 12f8c
		x"24690076", -- 12f90
		x"4e924e5e", -- 12f94
		x"2e9f4e75", -- 12f98
		x"4e750103", -- 12f9c
		x"01000800", -- 12fa0
		x"007d003e", -- 12fa4
		x"00a8005d", -- 12fa8
		x"0000007d", -- 12fac
		x"00000000", -- 12fb0
		x"00004e56", -- 12fb4
		x"fffc202e", -- 12fb8
		x"0008e580", -- 12fbc
		x"2d40fffc", -- 12fc0
		x"2f2efffc", -- 12fc4
		x"2f3c0000", -- 12fc8
		x"007d4eb9", -- 12fcc
		x"000081ac", -- 12fd0
		x"202efffc", -- 12fd4
		x"d09f2f00", -- 12fd8
		x"2f3c0000", -- 12fdc
		x"007d4eb9", -- 12fe0
		x"000081a8", -- 12fe4
		x"55972d5f", -- 12fe8
		x"000c4e5e", -- 12fec
		x"2e9f4e75", -- 12ff0
		x"00004e56", -- 12ff4
		x"fffc206e", -- 12ff8
		x"000c2068", -- 12ffc
		x"00482d68", -- 13000
		x"0044fffc", -- 13004
		x"206efffc", -- 13008
		x"117cff00", -- 1300c
		x"00111168", -- 13010
		x"00090009", -- 13014
		x"08e80007", -- 13018
		x"00112f3c", -- 1301c
		x"000f4240", -- 13020
		x"4eb90001", -- 13024
		x"4b16206e", -- 13028
		x"fffc4a28", -- 1302c
		x"000956c0", -- 13030
		x"66000012", -- 13034
		x"558f4eb9", -- 13038
		x"00014b30", -- 1303c
		x"101f6600", -- 13040
		x"000460e2", -- 13044
		x"206efffc", -- 13048
		x"08280005", -- 1304c
		x"000956c0", -- 13050
		x"44004a00", -- 13054
		x"67000010", -- 13058
		x"226e0008", -- 1305c
		x"22bc0000", -- 13060
		x"00036000", -- 13064
		x"001a2f2e", -- 13068
		x"000c3f3c", -- 1306c
		x"000e4eb9", -- 13070
		x"00011880", -- 13074
		x"206e0008", -- 13078
		x"20bc0000", -- 1307c
		x"0001206e", -- 13080
		x"fffc08a8", -- 13084
		x"00070011", -- 13088
		x"11680009", -- 1308c
		x"00094e5e", -- 13090
		x"205f504f", -- 13094
		x"4ed00000", -- 13098
		x"4e56fff0", -- 1309c
		x"2d6e000c", -- 130a0
		x"fffc206e", -- 130a4
		x"fffc2d68", -- 130a8
		x"0048fff8", -- 130ac
		x"226efff8", -- 130b0
		x"2d690040", -- 130b4
		x"fff42d69", -- 130b8
		x"0044fff0", -- 130bc
		x"4a280052", -- 130c0
		x"66000092", -- 130c4
		x"246e0008", -- 130c8
		x"24bc0000", -- 130cc
		x"0002117c", -- 130d0
		x"00010052", -- 130d4
		x"317c0014", -- 130d8
		x"0054246e", -- 130dc
		x"fff0156a", -- 130e0
		x"00090009", -- 130e4
		x"157c0000", -- 130e8
		x"0011598f", -- 130ec
		x"7000102a", -- 130f0
		x"00012f00", -- 130f4
		x"598f2f3c", -- 130f8
		x"00000001", -- 130fc
		x"30280002", -- 13100
		x"48c02f00", -- 13104
		x"4eb90001", -- 13108
		x"4b5a4eb9", -- 1310c
		x"00014b46", -- 13110
		x"201f206e", -- 13114
		x"fff01140", -- 13118
		x"00170228", -- 1311c
		x"001f0005", -- 13120
		x"7003eb88", -- 13124
		x"81280005", -- 13128
		x"42280019", -- 1312c
		x"117c0020", -- 13130
		x"001b117c", -- 13134
		x"0004001d", -- 13138
		x"0228001f", -- 1313c
		x"00057001", -- 13140
		x"eb888128", -- 13144
		x"0005226e", -- 13148
		x"fff408a9", -- 1314c
		x"00070003", -- 13150
		x"60000200", -- 13154
		x"206efffc", -- 13158
		x"42280052", -- 1315c
		x"226efff4", -- 13160
		x"08a90007", -- 13164
		x"0003246e", -- 13168
		x"fff0022a", -- 1316c
		x"ff1f0005", -- 13170
		x"7002eb88", -- 13174
		x"812a0005", -- 13178
		x"4a280053", -- 1317c
		x"67000010", -- 13180
		x"266e0008", -- 13184
		x"26bc0000", -- 13188
		x"00016000", -- 1318c
		x"01bc206e", -- 13190
		x"fff00828", -- 13194
		x"00020009", -- 13198
		x"56c04400", -- 1319c
		x"4a006700", -- 131a0
		x"0058226e", -- 131a4
		x"fffc7001", -- 131a8
		x"b0690056", -- 131ac
		x"66000034", -- 131b0
		x"246e0008", -- 131b4
		x"24bc0000", -- 131b8
		x"00012f2e", -- 131bc
		x"000c3f3c", -- 131c0
		x"00064eb9", -- 131c4
		x"00011880", -- 131c8
		x"206efff8", -- 131cc
		x"226efffc", -- 131d0
		x"30290002", -- 131d4
		x"48c0e580", -- 131d8
		x"31bc0001", -- 131dc
		x"08206000", -- 131e0
		x"0014206e", -- 131e4
		x"fffc5268", -- 131e8
		x"0056226e", -- 131ec
		x"000822bc", -- 131f0
		x"00000004", -- 131f4
		x"60000152", -- 131f8
		x"206efff0", -- 131fc
		x"08280004", -- 13200
		x"000956c0", -- 13204
		x"44004a00", -- 13208
		x"6700013e", -- 1320c
		x"1028000d", -- 13210
		x"e8880280", -- 13214
		x"0000000f", -- 13218
		x"7208b280", -- 1321c
		x"670000b4", -- 13220
		x"1028000d", -- 13224
		x"e8880280", -- 13228
		x"0000000f", -- 1322c
		x"7209b280", -- 13230
		x"670000a0", -- 13234
		x"2f3c000f", -- 13238
		x"42404eb9", -- 1323c
		x"00014b16", -- 13240
		x"206efff0", -- 13244
		x"1028000d", -- 13248
		x"e8880280", -- 1324c
		x"0000000f", -- 13250
		x"7208b280", -- 13254
		x"57c06700", -- 13258
		x"00281028", -- 1325c
		x"000de888", -- 13260
		x"02800000", -- 13264
		x"000f7209", -- 13268
		x"b28057c0", -- 1326c
		x"67000012", -- 13270
		x"558f4eb9", -- 13274
		x"00014b30", -- 13278
		x"101f6600", -- 1327c
		x"000460c0", -- 13280
		x"206efff0", -- 13284
		x"1028000d", -- 13288
		x"e8880280", -- 1328c
		x"0000000f", -- 13290
		x"7208b280", -- 13294
		x"67000032", -- 13298
		x"1028000d", -- 1329c
		x"e8880280", -- 132a0
		x"0000000f", -- 132a4
		x"7209b280", -- 132a8
		x"6700001e", -- 132ac
		x"206e0008", -- 132b0
		x"20bc0000", -- 132b4
		x"00012f2e", -- 132b8
		x"000c3f3c", -- 132bc
		x"000e4eb9", -- 132c0
		x"00011880", -- 132c4
		x"60000008", -- 132c8
		x"206e0008", -- 132cc
		x"42906000", -- 132d0
		x"0008206e", -- 132d4
		x"00084290", -- 132d8
		x"206efff0", -- 132dc
		x"1028000b", -- 132e0
		x"02800000", -- 132e4
		x"00077206", -- 132e8
		x"b2806700", -- 132ec
		x"005c1028", -- 132f0
		x"000b0280", -- 132f4
		x"00000007", -- 132f8
		x"7202b280", -- 132fc
		x"6700004a", -- 13300
		x"2f3c000f", -- 13304
		x"42404eb9", -- 13308
		x"00014b16", -- 1330c
		x"206efff0", -- 13310
		x"1028000b", -- 13314
		x"02800000", -- 13318
		x"00077206", -- 1331c
		x"b28057c0", -- 13320
		x"67000026", -- 13324
		x"1028000b", -- 13328
		x"02800000", -- 1332c
		x"00077202", -- 13330
		x"b28057c0", -- 13334
		x"67000012", -- 13338
		x"558f4eb9", -- 1333c
		x"00014b30", -- 13340
		x"101f6600", -- 13344
		x"000460c4", -- 13348
		x"206efff0", -- 1334c
		x"11680009", -- 13350
		x"00094e5e", -- 13354
		x"205f504f", -- 13358
		x"4ed00000", -- 1335c
		x"4e56ffee", -- 13360
		x"2d6e000c", -- 13364
		x"fff6206e", -- 13368
		x"fff62d68", -- 1336c
		x"0048fff2", -- 13370
		x"226efff2", -- 13374
		x"2d690044", -- 13378
		x"ffee7008", -- 1337c
		x"b0680004", -- 13380
		x"6f0000b8", -- 13384
		x"08ee0007", -- 13388
		x"fffe1028", -- 1338c
		x"00090840", -- 13390
		x"00000200", -- 13394
		x"000108ae", -- 13398
		x"0006fffe", -- 1339c
		x"ed88812e", -- 133a0
		x"fffe022e", -- 133a4
		x"ffc7fffe", -- 133a8
		x"7000e788", -- 133ac
		x"812efffe", -- 133b0
		x"022efff8", -- 133b4
		x"fffe3028", -- 133b8
		x"0004812e", -- 133bc
		x"fffe7000", -- 133c0
		x"102efffe", -- 133c4
		x"3d40fffc", -- 133c8
		x"30280002", -- 133cc
		x"48c0e580", -- 133d0
		x"4a710820", -- 133d4
		x"57c00200", -- 133d8
		x"08011d40", -- 133dc
		x"fffb558f", -- 133e0
		x"2f2e000c", -- 133e4
		x"486efffc", -- 133e8
		x"3f3c0006", -- 133ec
		x"1f2efffb", -- 133f0
		x"42274eb9", -- 133f4
		x"00012454", -- 133f8
		x"4a1f6700", -- 133fc
		x"00224a2e", -- 13400
		x"fffb6700", -- 13404
		x"0010206e", -- 13408
		x"000820bc", -- 1340c
		x"00000013", -- 13410
		x"60000008", -- 13414
		x"206e0008", -- 13418
		x"42906000", -- 1341c
		x"001a2f2e", -- 13420
		x"000c3f3c", -- 13424
		x"00074eb9", -- 13428
		x"00011880", -- 1342c
		x"206e0008", -- 13430
		x"20bc0000", -- 13434
		x"00016000", -- 13438
		x"001a2f2e", -- 1343c
		x"000c3f3c", -- 13440
		x"00054eb9", -- 13444
		x"00011880", -- 13448
		x"206e0008", -- 1344c
		x"20bc0000", -- 13450
		x"00014e5e", -- 13454
		x"205f504f", -- 13458
		x"4ed00000", -- 1345c
		x"4e56ffce", -- 13460
		x"2d6e000c", -- 13464
		x"ffe2206e", -- 13468
		x"ffe22d68", -- 1346c
		x"0048ffde", -- 13470
		x"226effde", -- 13474
		x"2d690040", -- 13478
		x"ffda2d69", -- 1347c
		x"0044ffd6", -- 13480
		x"30280002", -- 13484
		x"48c0e580", -- 13488
		x"45f10820", -- 1348c
		x"2d4affd2", -- 13490
		x"246e0008", -- 13494
		x"42922d7a", -- 13498
		x"fb02fffa", -- 1349c
		x"1d7afb00", -- 134a0
		x"fffe558f", -- 134a4
		x"2d40ffce", -- 134a8
		x"4eb90001", -- 134ac
		x"1a92202e", -- 134b0
		x"ffce101f", -- 134b4
		x"67000016", -- 134b8
		x"206effda", -- 134bc
		x"08280005", -- 134c0
		x"000156c1", -- 134c4
		x"44010841", -- 134c8
		x"00001001", -- 134cc
		x"02000001", -- 134d0
		x"72001200", -- 134d4
		x"2d41fff0", -- 134d8
		x"206effda", -- 134dc
		x"10280007", -- 134e0
		x"ea880280", -- 134e4
		x"00000003", -- 134e8
		x"e580222e", -- 134ec
		x"fff0d281", -- 134f0
		x"d28043fa", -- 134f4
		x"faac1d71", -- 134f8
		x"1801fffd", -- 134fc
		x"4a2efffd", -- 13500
		x"66000054", -- 13504
		x"226effd2", -- 13508
		x"32bc0001", -- 1350c
		x"3d7c0008", -- 13510
		x"ffee558f", -- 13514
		x"2f2e000c", -- 13518
		x"486effee", -- 1351c
		x"3f3c0006", -- 13520
		x"42274227", -- 13524
		x"4eb90001", -- 13528
		x"24544a1f", -- 1352c
		x"6600001e", -- 13530
		x"206e0008", -- 13534
		x"20bc0000", -- 13538
		x"00012f2e", -- 1353c
		x"000c3f3c", -- 13540
		x"00074eb9", -- 13544
		x"00011880", -- 13548
		x"60000008", -- 1354c
		x"206e0008", -- 13550
		x"42906000", -- 13554
		x"028e41ee", -- 13558
		x"fffa2d48", -- 1355c
		x"ffe62d7c", -- 13560
		x"00000005", -- 13564
		x"ffea7000", -- 13568
		x"206effe6", -- 1356c
		x"10103d40", -- 13570
		x"ffee206e", -- 13574
		x"ffd61028", -- 13578
		x"000b0280", -- 1357c
		x"00000007", -- 13580
		x"7206b280", -- 13584
		x"66000090", -- 13588
		x"4aaeffea", -- 1358c
		x"6f000088", -- 13590
		x"206e0008", -- 13594
		x"4a906600", -- 13598
		x"007e558f", -- 1359c
		x"2f2e000c", -- 135a0
		x"486effee", -- 135a4
		x"3f3c0006", -- 135a8
		x"7001b0ae", -- 135ac
		x"ffea5dc0", -- 135b0
		x"0200ff01", -- 135b4
		x"1f004227", -- 135b8
		x"4eb90001", -- 135bc
		x"24544a1f", -- 135c0
		x"6700001a", -- 135c4
		x"52aeffe6", -- 135c8
		x"7000206e", -- 135cc
		x"ffe61010", -- 135d0
		x"3d40ffee", -- 135d4
		x"53aeffea", -- 135d8
		x"60000038", -- 135dc
		x"206effd6", -- 135e0
		x"1028000b", -- 135e4
		x"02800000", -- 135e8
		x"00077206", -- 135ec
		x"b2806600", -- 135f0
		x"0022226e", -- 135f4
		x"ffd232bc", -- 135f8
		x"0001246e", -- 135fc
		x"000824bc", -- 13600
		x"00000001", -- 13604
		x"2f2e000c", -- 13608
		x"3f3c0007", -- 1360c
		x"4eb90001", -- 13610
		x"18806000", -- 13614
		x"ff5e206e", -- 13618
		x"00084a90", -- 1361c
		x"660001c4", -- 13620
		x"41eefff4", -- 13624
		x"2d48ffe6", -- 13628
		x"42aeffea", -- 1362c
		x"206effd6", -- 13630
		x"1028000b", -- 13634
		x"02800000", -- 13638
		x"00077207", -- 1363c
		x"b2806600", -- 13640
		x"0084226e", -- 13644
		x"00084a91", -- 13648
		x"6600007a", -- 1364c
		x"558f2f2e", -- 13650
		x"000c486e", -- 13654
		x"ffee3f3c", -- 13658
		x"00077004", -- 1365c
		x"b0aeffea", -- 13660
		x"5ec00200", -- 13664
		x"ff011f00", -- 13668
		x"42274eb9", -- 1366c
		x"00012454", -- 13670
		x"4a1f6700", -- 13674
		x"0016206e", -- 13678
		x"ffe610ae", -- 1367c
		x"ffef52ae", -- 13680
		x"ffe652ae", -- 13684
		x"ffea6000", -- 13688
		x"0038206e", -- 1368c
		x"ffd61028", -- 13690
		x"000b0280", -- 13694
		x"00000007", -- 13698
		x"7207b280", -- 1369c
		x"66000022", -- 136a0
		x"226effd2", -- 136a4
		x"32bc0001", -- 136a8
		x"246e0008", -- 136ac
		x"24bc0000", -- 136b0
		x"00012f2e", -- 136b4
		x"000c3f3c", -- 136b8
		x"00074eb9", -- 136bc
		x"00011880", -- 136c0
		x"6000ff6a", -- 136c4
		x"206e0008", -- 136c8
		x"4a906600", -- 136cc
		x"01064aae", -- 136d0
		x"ffea6f00", -- 136d4
		x"00fe7001", -- 136d8
		x"b0aeffea", -- 136dc
		x"66000018", -- 136e0
		x"7007b02e", -- 136e4
		x"fff46600", -- 136e8
		x"000e206e", -- 136ec
		x"ffd230bc", -- 136f0
		x"00016000", -- 136f4
		x"00da7005", -- 136f8
		x"b0aeffea", -- 136fc
		x"660000ba", -- 13700
		x"7001b02e", -- 13704
		x"fff46600", -- 13708
		x"00b07001", -- 1370c
		x"b02efff6", -- 13710
		x"660000a6", -- 13714
		x"4a2efff8", -- 13718
		x"6600000e", -- 1371c
		x"206effd2", -- 13720
		x"30bc0001", -- 13724
		x"6000008e", -- 13728
		x"598f7000", -- 1372c
		x"102efff7", -- 13730
		x"2f004eba", -- 13734
		x"f87e2d5f", -- 13738
		x"ffea102e", -- 1373c
		x"fff8b02e", -- 13740
		x"fffe6200", -- 13744
		x"005a102e", -- 13748
		x"fff7b02e", -- 1374c
		x"fffd6500", -- 13750
		x"004e7004", -- 13754
		x"b0aeffea", -- 13758
		x"6f000044", -- 1375c
		x"206effd2", -- 13760
		x"30bc0002", -- 13764
		x"08e80007", -- 13768
		x"0003102e", -- 1376c
		x"fffe0200", -- 13770
		x"ff070228", -- 13774
		x"ff8f0003", -- 13778
		x"e9888128", -- 1377c
		x"00030228", -- 13780
		x"00f30003", -- 13784
		x"202effea", -- 13788
		x"e5888128", -- 1378c
		x"00030228", -- 13790
		x"00fc0003", -- 13794
		x"70008128", -- 13798
		x"00036000", -- 1379c
		x"0018206e", -- 137a0
		x"ffd230bc", -- 137a4
		x"00012f2e", -- 137a8
		x"000c2f2e", -- 137ac
		x"00084eb9", -- 137b0
		x"00013c50", -- 137b4
		x"60000018", -- 137b8
		x"206effd2", -- 137bc
		x"30bc0001", -- 137c0
		x"2f2e000c", -- 137c4
		x"2f2e0008", -- 137c8
		x"4eb90001", -- 137cc
		x"3c506000", -- 137d0
		x"00124aae", -- 137d4
		x"ffea6600", -- 137d8
		x"000a206e", -- 137dc
		x"ffd230bc", -- 137e0
		x"00014e5e", -- 137e4
		x"205f504f", -- 137e8
		x"4ed00000", -- 137ec
		x"4e56ffcc", -- 137f0
		x"2d6e000c", -- 137f4
		x"ffe4206e", -- 137f8
		x"ffe443e8", -- 137fc
		x"00442d49", -- 13800
		x"ffe0226e", -- 13804
		x"ffe02d69", -- 13808
		x"0004ffdc", -- 1380c
		x"246effdc", -- 13810
		x"2d6a0040", -- 13814
		x"ffd82d6a", -- 13818
		x"0044ffd4", -- 1381c
		x"30280002", -- 13820
		x"48c0e580", -- 13824
		x"47f20820", -- 13828
		x"2d4bffd0", -- 1382c
		x"266effd0", -- 13830
		x"4253286e", -- 13834
		x"00084294", -- 13838
		x"2d7af760", -- 1383c
		x"fffa1d7a", -- 13840
		x"f75efffe", -- 13844
		x"558f2d40", -- 13848
		x"ffcc4eb9", -- 1384c
		x"00011a92", -- 13850
		x"202effcc", -- 13854
		x"101f6700", -- 13858
		x"0016206e", -- 1385c
		x"ffd80828", -- 13860
		x"00050001", -- 13864
		x"56c14401", -- 13868
		x"08410000", -- 1386c
		x"10010200", -- 13870
		x"00017200", -- 13874
		x"12002d41", -- 13878
		x"fff64a2e", -- 1387c
		x"fffd6600", -- 13880
		x"001c206e", -- 13884
		x"ffd030bc", -- 13888
		x"00012f2e", -- 1388c
		x"000c2f2e", -- 13890
		x"00084eb9", -- 13894
		x"00013c50", -- 13898
		x"600001aa", -- 1389c
		x"206effe0", -- 138a0
		x"4a68002e", -- 138a4
		x"6600001c", -- 138a8
		x"226effd0", -- 138ac
		x"32bc0001", -- 138b0
		x"2f2e000c", -- 138b4
		x"2f2e0008", -- 138b8
		x"4eb90001", -- 138bc
		x"3c506000", -- 138c0
		x"001a206e", -- 138c4
		x"ffe07000", -- 138c8
		x"102efffe", -- 138cc
		x"b068002e", -- 138d0
		x"6f000008", -- 138d4
		x"1d68002f", -- 138d8
		x"fffe206e", -- 138dc
		x"ffe07000", -- 138e0
		x"102efffd", -- 138e4
		x"b0680030", -- 138e8
		x"6c000046", -- 138ec
		x"598f3028", -- 138f0
		x"003048c0", -- 138f4
		x"2f004eba", -- 138f8
		x"f6ba2d5f", -- 138fc
		x"ffec7004", -- 13900
		x"b0aeffec", -- 13904
		x"6f000010", -- 13908
		x"206effe0", -- 1390c
		x"1d680031", -- 13910
		x"fffd6000", -- 13914
		x"0018206e", -- 13918
		x"ffd030bc", -- 1391c
		x"00012f2e", -- 13920
		x"000c2f2e", -- 13924
		x"00084eb9", -- 13928
		x"00013c50", -- 1392c
		x"60000014", -- 13930
		x"598f7000", -- 13934
		x"102efffd", -- 13938
		x"2f004eba", -- 1393c
		x"f6762d5f", -- 13940
		x"ffec206e", -- 13944
		x"ffd04a50", -- 13948
		x"660000fa", -- 1394c
		x"226e0008", -- 13950
		x"429143ee", -- 13954
		x"fffa2d49", -- 13958
		x"ffe82d7c", -- 1395c
		x"00000005", -- 13960
		x"fff07000", -- 13964
		x"226effe8", -- 13968
		x"10113d40", -- 1396c
		x"fff4206e", -- 13970
		x"ffd41028", -- 13974
		x"000b0280", -- 13978
		x"00000007", -- 1397c
		x"7206b280", -- 13980
		x"6600007a", -- 13984
		x"4aaefff0", -- 13988
		x"6f000072", -- 1398c
		x"206e0008", -- 13990
		x"4a906600", -- 13994
		x"0068558f", -- 13998
		x"2f2e000c", -- 1399c
		x"486efff4", -- 139a0
		x"3f3c0006", -- 139a4
		x"7001b0ae", -- 139a8
		x"fff05dc0", -- 139ac
		x"0200ff01", -- 139b0
		x"1f004227", -- 139b4
		x"4eb90001", -- 139b8
		x"24544a1f", -- 139bc
		x"6700001a", -- 139c0
		x"52aeffe8", -- 139c4
		x"7000206e", -- 139c8
		x"ffe81010", -- 139cc
		x"3d40fff4", -- 139d0
		x"53aefff0", -- 139d4
		x"60000022", -- 139d8
		x"206effd0", -- 139dc
		x"30bc0001", -- 139e0
		x"226e0008", -- 139e4
		x"22bc0000", -- 139e8
		x"00012f2e", -- 139ec
		x"000c3f3c", -- 139f0
		x"00074eb9", -- 139f4
		x"00011880", -- 139f8
		x"6000ff74", -- 139fc
		x"206e0008", -- 13a00
		x"4a906600", -- 13a04
		x"0040206e", -- 13a08
		x"ffd030bc", -- 13a0c
		x"000208e8", -- 13a10
		x"00070003", -- 13a14
		x"102efffe", -- 13a18
		x"0200ff07", -- 13a1c
		x"0228ff8f", -- 13a20
		x"0003e988", -- 13a24
		x"81280003", -- 13a28
		x"022800f3", -- 13a2c
		x"0003202e", -- 13a30
		x"ffece588", -- 13a34
		x"81280003", -- 13a38
		x"022800fc", -- 13a3c
		x"00037000", -- 13a40
		x"81280003", -- 13a44
		x"4e5e205f", -- 13a48
		x"504f4ed0", -- 13a4c
		x"0000000e", -- 13a50
		x"00000001", -- 13a54
		x"0000000b", -- 13a58
		x"0000000c", -- 13a5c
		x"0000000d", -- 13a60
		x"00000001", -- 13a64
		x"00000001", -- 13a68
		x"00000001", -- 13a6c
		x"00000001", -- 13a70
		x"00000001", -- 13a74
		x"00000011", -- 13a78
		x"00000012", -- 13a7c
		x"00000001", -- 13a80
		x"00004e56", -- 13a84
		x"ffec206e", -- 13a88
		x"000c41e8", -- 13a8c
		x"00442d48", -- 13a90
		x"fff0206e", -- 13a94
		x"fff02268", -- 13a98
		x"00042d69", -- 13a9c
		x"0044ffec", -- 13aa0
		x"226e0008", -- 13aa4
		x"429142ae", -- 13aa8
		x"fff4206e", -- 13aac
		x"ffec1028", -- 13ab0
		x"000b0280", -- 13ab4
		x"00000007", -- 13ab8
		x"7207b280", -- 13abc
		x"660000a4", -- 13ac0
		x"226e0008", -- 13ac4
		x"4a916600", -- 13ac8
		x"009a558f", -- 13acc
		x"2f2e000c", -- 13ad0
		x"486efff8", -- 13ad4
		x"3f3c0007", -- 13ad8
		x"7004b0ae", -- 13adc
		x"fff45ec0", -- 13ae0
		x"0200ff01", -- 13ae4
		x"1f007204", -- 13ae8
		x"b2aefff4", -- 13aec
		x"57c11001", -- 13af0
		x"6700001a", -- 13af4
		x"7201b22e", -- 13af8
		x"fffa57c1", -- 13afc
		x"10016700", -- 13b00
		x"000c7201", -- 13b04
		x"b22efffc", -- 13b08
		x"57c11001", -- 13b0c
		x"0200ff01", -- 13b10
		x"1f004eb9", -- 13b14
		x"00012454", -- 13b18
		x"4a1f6700", -- 13b1c
		x"001452ae", -- 13b20
		x"fff4202e", -- 13b24
		x"fff41dae", -- 13b28
		x"fff908f9", -- 13b2c
		x"60000030", -- 13b30
		x"206effec", -- 13b34
		x"1028000b", -- 13b38
		x"02800000", -- 13b3c
		x"00077207", -- 13b40
		x"b2806600", -- 13b44
		x"001a226e", -- 13b48
		x"000822bc", -- 13b4c
		x"00000001", -- 13b50
		x"2f2e000c", -- 13b54
		x"3f3c0007", -- 13b58
		x"4eb90001", -- 13b5c
		x"18806000", -- 13b60
		x"ff4a7000", -- 13b64
		x"102efffa", -- 13b68
		x"3d40fff8", -- 13b6c
		x"7001b0ae", -- 13b70
		x"fff46600", -- 13b74
		x"0050302e", -- 13b78
		x"fff86c04", -- 13b7c
		x"d07c007f", -- 13b80
		x"ee406700", -- 13b84
		x"0010206e", -- 13b88
		x"000820bc", -- 13b8c
		x"00000010", -- 13b90
		x"6000002e", -- 13b94
		x"700cb06e", -- 13b98
		x"fff86c00", -- 13b9c
		x"0010206e", -- 13ba0
		x"000820bc", -- 13ba4
		x"00000001", -- 13ba8
		x"60000016", -- 13bac
		x"302efff8", -- 13bb0
		x"48c0e580", -- 13bb4
		x"206e0008", -- 13bb8
		x"43fafe92", -- 13bbc
		x"20b10800", -- 13bc0
		x"60000066", -- 13bc4
		x"7001b06e", -- 13bc8
		x"fff86600", -- 13bcc
		x"00527005", -- 13bd0
		x"b0aefff4", -- 13bd4
		x"66000048", -- 13bd8
		x"7001b02e", -- 13bdc
		x"fffc6600", -- 13be0
		x"003e206e", -- 13be4
		x"ffec1028", -- 13be8
		x"000b0280", -- 13bec
		x"00000007", -- 13bf0
		x"7206b280", -- 13bf4
		x"66000028", -- 13bf8
		x"206e0008", -- 13bfc
		x"20bc0000", -- 13c00
		x"000a206e", -- 13c04
		x"fff07000", -- 13c08
		x"102efffd", -- 13c0c
		x"31400030", -- 13c10
		x"7000102e", -- 13c14
		x"fffe3140", -- 13c18
		x"002e6000", -- 13c1c
		x"000c206e", -- 13c20
		x"000820bc", -- 13c24
		x"00000001", -- 13c28
		x"206e0008", -- 13c2c
		x"7001b090", -- 13c30
		x"66000010", -- 13c34
		x"2f2e000c", -- 13c38
		x"3f3c000d", -- 13c3c
		x"4eb90001", -- 13c40
		x"18804e5e", -- 13c44
		x"205f504f", -- 13c48
		x"4ed00000", -- 13c4c
		x"4e56fffe", -- 13c50
		x"2f2e000c", -- 13c54
		x"2f2e0008", -- 13c58
		x"4eb90001", -- 13c5c
		x"207a206e", -- 13c60
		x"00087006", -- 13c64
		x"b0906600", -- 13c68
		x"00483d7c", -- 13c6c
		x"0007fffe", -- 13c70
		x"558f2f2e", -- 13c74
		x"000c486e", -- 13c78
		x"fffe3f3c", -- 13c7c
		x"00064227", -- 13c80
		x"42274eb9", -- 13c84
		x"00012454", -- 13c88
		x"4a1f6700", -- 13c8c
		x"000c206e", -- 13c90
		x"00084290", -- 13c94
		x"6000001a", -- 13c98
		x"206e0008", -- 13c9c
		x"20bc0000", -- 13ca0
		x"00012f2e", -- 13ca4
		x"000c3f3c", -- 13ca8
		x"00074eb9", -- 13cac
		x"00011880", -- 13cb0
		x"4e5e205f", -- 13cb4
		x"504f4ed0", -- 13cb8
		x"00004e56", -- 13cbc
		x"ffee206e", -- 13cc0
		x"00084290", -- 13cc4
		x"2d6e000c", -- 13cc8
		x"fffa206e", -- 13ccc
		x"fffa43e8", -- 13cd0
		x"00582d49", -- 13cd4
		x"fff62d68", -- 13cd8
		x"0048fff2", -- 13cdc
		x"226efff2", -- 13ce0
		x"30280002", -- 13ce4
		x"48c0e580", -- 13ce8
		x"45f10820", -- 13cec
		x"2d4affee", -- 13cf0
		x"24690044", -- 13cf4
		x"266efff6", -- 13cf8
		x"102a000b", -- 13cfc
		x"02800000", -- 13d00
		x"00073680", -- 13d04
		x"426b0002", -- 13d08
		x"30136d00", -- 13d0c
		x"0098b07c", -- 13d10
		x"00026e00", -- 13d14
		x"0090e340", -- 13d18
		x"323b0006", -- 13d1c
		x"4efb1002", -- 13d20
		x"00480066", -- 13d24
		x"00062768", -- 13d28
		x"000a0010", -- 13d2c
		x"3028000e", -- 13d30
		x"48c02740", -- 13d34
		x"0014422b", -- 13d38
		x"0018246e", -- 13d3c
		x"ffee7002", -- 13d40
		x"b0526600", -- 13d44
		x"000c1d6a", -- 13d48
		x"0003ffff", -- 13d4c
		x"60000008", -- 13d50
		x"1d7c0000", -- 13d54
		x"ffff206e", -- 13d58
		x"fff22268", -- 13d5c
		x"0044136e", -- 13d60
		x"ffff0007", -- 13d64
		x"60000056", -- 13d68
		x"206efffa", -- 13d6c
		x"226efff6", -- 13d70
		x"4ca81c01", -- 13d74
		x"001a48a9", -- 13d78
		x"1c010010", -- 13d7c
		x"13680022", -- 13d80
		x"00186000", -- 13d84
		x"0038206e", -- 13d88
		x"fffa226e", -- 13d8c
		x"fff64ca8", -- 13d90
		x"1c010010", -- 13d94
		x"48a91c01", -- 13d98
		x"00101368", -- 13d9c
		x"00180018", -- 13da0
		x"6000001a", -- 13da4
		x"2f2e000c", -- 13da8
		x"3f3c000b", -- 13dac
		x"4eb90001", -- 13db0
		x"1880206e", -- 13db4
		x"000820bc", -- 13db8
		x"00000001", -- 13dbc
		x"206e0008", -- 13dc0
		x"4a906600", -- 13dc4
		x"0012206e", -- 13dc8
		x"fff62168", -- 13dcc
		x"00100004", -- 13dd0
		x"21680014", -- 13dd4
		x"00084e5e", -- 13dd8
		x"205f504f", -- 13ddc
		x"4ed00000", -- 13de0
		x"4e560000", -- 13de4
		x"206e0008", -- 13de8
		x"42904e5e", -- 13dec
		x"205f504f", -- 13df0
		x"4ed00000", -- 13df4
		x"4e56ffec", -- 13df8
		x"2d6e000c", -- 13dfc
		x"fffc206e", -- 13e00
		x"fffc43e8", -- 13e04
		x"00442d49", -- 13e08
		x"fff8226e", -- 13e0c
		x"fff845e9", -- 13e10
		x"00142d4a", -- 13e14
		x"fff42d69", -- 13e18
		x"0004fff0", -- 13e1c
		x"246efff0", -- 13e20
		x"2d6a0044", -- 13e24
		x"ffec266e", -- 13e28
		x"00084293", -- 13e2c
		x"4a29000e", -- 13e30
		x"66000092", -- 13e34
		x"4a29002c", -- 13e38
		x"67000026", -- 13e3c
		x"598f3f10", -- 13e40
		x"4eb90001", -- 13e44
		x"1afa206e", -- 13e48
		x"fff0215f", -- 13e4c
		x"004e70ff", -- 13e50
		x"b0a8004e", -- 13e54
		x"6600000a", -- 13e58
		x"226efff4", -- 13e5c
		x"42290018", -- 13e60
		x"206efff8", -- 13e64
		x"4a28002c", -- 13e68
		x"6700003a", -- 13e6c
		x"226efff0", -- 13e70
		x"137cff01", -- 13e74
		x"004c558f", -- 13e78
		x"2f2e000c", -- 13e7c
		x"4eb90001", -- 13e80
		x"26f64a1f", -- 13e84
		x"66000010", -- 13e88
		x"206e0008", -- 13e8c
		x"20bc0000", -- 13e90
		x"00016000", -- 13e94
		x"000c206e", -- 13e98
		x"000820bc", -- 13e9c
		x"00000002", -- 13ea0
		x"6000001e", -- 13ea4
		x"558f2f2e", -- 13ea8
		x"000c4eb9", -- 13eac
		x"00012ae2", -- 13eb0
		x"4a1f6600", -- 13eb4
		x"000c206e", -- 13eb8
		x"000820bc", -- 13ebc
		x"00000001", -- 13ec0
		x"60000064", -- 13ec4
		x"558f2f2e", -- 13ec8
		x"000c2f2e", -- 13ecc
		x"00084eb9", -- 13ed0
		x"000128e2", -- 13ed4
		x"4a1f6600", -- 13ed8
		x"003a206e", -- 13edc
		x"fff0117c", -- 13ee0
		x"ff01004c", -- 13ee4
		x"558f2f2e", -- 13ee8
		x"000c4eb9", -- 13eec
		x"000126f6", -- 13ef0
		x"4a1f6600", -- 13ef4
		x"0010206e", -- 13ef8
		x"000820bc", -- 13efc
		x"00000001", -- 13f00
		x"6000000c", -- 13f04
		x"206e0008", -- 13f08
		x"20bc0000", -- 13f0c
		x"00026000", -- 13f10
		x"0016206e", -- 13f14
		x"fffc3f10", -- 13f18
		x"4eb90001", -- 13f1c
		x"1f28206e", -- 13f20
		x"fff04228", -- 13f24
		x"004c206e", -- 13f28
		x"00084a90", -- 13f2c
		x"6600007c", -- 13f30
		x"206efff4", -- 13f34
		x"226effec", -- 13f38
		x"1029000b", -- 13f3c
		x"02800000", -- 13f40
		x"00073210", -- 13f44
		x"48c1b280", -- 13f48
		x"66000060", -- 13f4c
		x"206efff4", -- 13f50
		x"226effec", -- 13f54
		x"1029000b", -- 13f58
		x"02800000", -- 13f5c
		x"00073210", -- 13f60
		x"48c1b280", -- 13f64
		x"56c06600", -- 13f68
		x"000e4a29", -- 13f6c
		x"000956c0", -- 13f70
		x"66000004", -- 13f74
		x"60d6206e", -- 13f78
		x"fff4226e", -- 13f7c
		x"ffec1029", -- 13f80
		x"000b0280", -- 13f84
		x"00000007", -- 13f88
		x"321048c1", -- 13f8c
		x"b2806600", -- 13f90
		x"001a246e", -- 13f94
		x"000824bc", -- 13f98
		x"00000001", -- 13f9c
		x"2f2e000c", -- 13fa0
		x"3f3c0008", -- 13fa4
		x"4eb90001", -- 13fa8
		x"18804e5e", -- 13fac
		x"205f504f", -- 13fb0
		x"4ed00000", -- 13fb4
		x"4e56fffa", -- 13fb8
		x"206e000c", -- 13fbc
		x"41e80058", -- 13fc0
		x"2d48fffa", -- 13fc4
		x"206efffa", -- 13fc8
		x"52680002", -- 13fcc
		x"7002b068", -- 13fd0
		x"00026c00", -- 13fd4
		x"001e226e", -- 13fd8
		x"000822bc", -- 13fdc
		x"00000001", -- 13fe0
		x"2f2e000c", -- 13fe4
		x"3f3c0009", -- 13fe8
		x"4eb90001", -- 13fec
		x"18806000", -- 13ff0
		x"00483d7c", -- 13ff4
		x"0005fffe", -- 13ff8
		x"558f2f2e", -- 13ffc
		x"000c486e", -- 14000
		x"fffe3f3c", -- 14004
		x"00064227", -- 14008
		x"42274eb9", -- 1400c
		x"00012454", -- 14010
		x"4a1f6700", -- 14014
		x"000c206e", -- 14018
		x"00084290", -- 1401c
		x"6000001a", -- 14020
		x"206e0008", -- 14024
		x"20bc0000", -- 14028
		x"00012f2e", -- 1402c
		x"000c3f3c", -- 14030
		x"00084eb9", -- 14034
		x"00011880", -- 14038
		x"4e5e205f", -- 1403c
		x"504f4ed0", -- 14040
		x"00004e56", -- 14044
		x"ffee206e", -- 14048
		x"000c41e8", -- 1404c
		x"00442d48", -- 14050
		x"fff2206e", -- 14054
		x"fff243e8", -- 14058
		x"00142d49", -- 1405c
		x"ffee4a68", -- 14060
		x"003a6600", -- 14064
		x"0016226e", -- 14068
		x"ffee2369", -- 1406c
		x"00100004", -- 14070
		x"23690014", -- 14074
		x"00086000", -- 14078
		x"0160206e", -- 1407c
		x"ffee2028", -- 14080
		x"000890a8", -- 14084
		x"00142d40", -- 14088
		x"fffc3d7c", -- 1408c
		x"0001fffa", -- 14090
		x"426efff6", -- 14094
		x"526efff6", -- 14098
		x"206efff2", -- 1409c
		x"302efff6", -- 140a0
		x"48c0d080", -- 140a4
		x"4a700838", -- 140a8
		x"6f00007a", -- 140ac
		x"302efff6", -- 140b0
		x"48c0d080", -- 140b4
		x"30300838", -- 140b8
		x"48c0b0ae", -- 140bc
		x"fffc6d00", -- 140c0
		x"000c3d6e", -- 140c4
		x"fffefff8", -- 140c8
		x"60000014", -- 140cc
		x"206efff2", -- 140d0
		x"302efff6", -- 140d4
		x"48c0d080", -- 140d8
		x"3d700838", -- 140dc
		x"fff8206e", -- 140e0
		x"ffee302e", -- 140e4
		x"fff848c0", -- 140e8
		x"d1a80004", -- 140ec
		x"302efff8", -- 140f0
		x"48c091a8", -- 140f4
		x"0008302e", -- 140f8
		x"fff848c0", -- 140fc
		x"91aefffc", -- 14100
		x"226efff2", -- 14104
		x"302efff6", -- 14108
		x"48c0d080", -- 1410c
		x"30310838", -- 14110
		x"906efff8", -- 14114
		x"322efffa", -- 14118
		x"48c1d281", -- 1411c
		x"33801838", -- 14120
		x"6000007a", -- 14124
		x"206efff2", -- 14128
		x"302efff6", -- 1412c
		x"48c0d080", -- 14130
		x"4a700838", -- 14134
		x"6c000066", -- 14138
		x"302efff6", -- 1413c
		x"48c0d080", -- 14140
		x"30300838", -- 14144
		x"48c06c02", -- 14148
		x"4480b0ae", -- 1414c
		x"fffc6d00", -- 14150
		x"000c3d6e", -- 14154
		x"fffefff8", -- 14158
		x"60000018", -- 1415c
		x"206efff2", -- 14160
		x"302efff6", -- 14164
		x"48c0d080", -- 14168
		x"30300838", -- 1416c
		x"44403d40", -- 14170
		x"fff8302e", -- 14174
		x"fff848c0", -- 14178
		x"91aefffc", -- 1417c
		x"206efff2", -- 14180
		x"302efff6", -- 14184
		x"48c0d080", -- 14188
		x"30300838", -- 1418c
		x"d06efff8", -- 14190
		x"322efffa", -- 14194
		x"48c1d281", -- 14198
		x"31801838", -- 1419c
		x"206efff2", -- 141a0
		x"302efff6", -- 141a4
		x"48c0d080", -- 141a8
		x"4a700838", -- 141ac
		x"67000006", -- 141b0
		x"526efffa", -- 141b4
		x"0c6e0003", -- 141b8
		x"fff66d00", -- 141bc
		x"fed87004", -- 141c0
		x"b06efffa", -- 141c4
		x"6f000012", -- 141c8
		x"206efff2", -- 141cc
		x"302efffa", -- 141d0
		x"48c0d080", -- 141d4
		x"42700838", -- 141d8
		x"206e0008", -- 141dc
		x"42904e5e", -- 141e0
		x"205f504f", -- 141e4
		x"4ed00000", -- 141e8
		x"4e560000", -- 141ec
		x"206e000c", -- 141f0
		x"317c0002", -- 141f4
		x"002c206e", -- 141f8
		x"00084290", -- 141fc
		x"4e5e205f", -- 14200
		x"504f4ed0", -- 14204
		x"00004e56", -- 14208
		x"fffc206e", -- 1420c
		x"000c41e8", -- 14210
		x"00582d48", -- 14214
		x"fffc206e", -- 14218
		x"fffc2168", -- 1421c
		x"00040010", -- 14220
		x"21680008", -- 14224
		x"0014206e", -- 14228
		x"00084290", -- 1422c
		x"4e5e205f", -- 14230
		x"504f4ed0", -- 14234
		x"00004e56", -- 14238
		x"fff82f2e", -- 1423c
		x"000c2f2e", -- 14240
		x"00084eb9", -- 14244
		x"00011f7c", -- 14248
		x"206e000c", -- 1424c
		x"41e80058", -- 14250
		x"2d48fffc", -- 14254
		x"206e000c", -- 14258
		x"20680048", -- 1425c
		x"2d680044", -- 14260
		x"fff8206e", -- 14264
		x"00087007", -- 14268
		x"b0906600", -- 1426c
		x"001c206e", -- 14270
		x"fffc7002", -- 14274
		x"b0506600", -- 14278
		x"0010206e", -- 1427c
		x"000820bc", -- 14280
		x"00000014", -- 14284
		x"60000050", -- 14288
		x"206e0008", -- 1428c
		x"7008b090", -- 14290
		x"66000044", -- 14294
		x"206efff8", -- 14298
		x"08280000", -- 1429c
		x"000b56c0", -- 142a0
		x"44004a00", -- 142a4
		x"6700001c", -- 142a8
		x"226efffc", -- 142ac
		x"7001b051", -- 142b0
		x"6600000c", -- 142b4
		x"246e0008", -- 142b8
		x"24bc0000", -- 142bc
		x"00146000", -- 142c0
		x"0016206e", -- 142c4
		x"fffc4a50", -- 142c8
		x"6600000c", -- 142cc
		x"226e0008", -- 142d0
		x"22bc0000", -- 142d4
		x"00144e5e", -- 142d8
		x"205f504f", -- 142dc
		x"4ed00000", -- 142e0
		x"4e56ffe4", -- 142e4
		x"2d6e000c", -- 142e8
		x"fff8206e", -- 142ec
		x"fff843e8", -- 142f0
		x"00442d49", -- 142f4
		x"fff4226e", -- 142f8
		x"fff42d69", -- 142fc
		x"0004fff0", -- 14300
		x"246efff0", -- 14304
		x"2d6a0040", -- 14308
		x"ffec2d6a", -- 1430c
		x"0044ffe8", -- 14310
		x"30280002", -- 14314
		x"48c0e580", -- 14318
		x"47f20820", -- 1431c
		x"2d4bffe4", -- 14320
		x"4a29000e", -- 14324
		x"66000036", -- 14328
		x"266e0008", -- 1432c
		x"26bc0000", -- 14330
		x"0002137c", -- 14334
		x"0001000e", -- 14338
		x"337c0040", -- 1433c
		x"0010266e", -- 14340
		x"ffe8176b", -- 14344
		x"00090009", -- 14348
		x"08eb0001", -- 1434c
		x"0003286e", -- 14350
		x"ffec08ac", -- 14354
		x"00070003", -- 14358
		x"600000f4", -- 1435c
		x"206effec", -- 14360
		x"08a80007", -- 14364
		x"0003226e", -- 14368
		x"ffe808a9", -- 1436c
		x"00010003", -- 14370
		x"246efff4", -- 14374
		x"422a000e", -- 14378
		x"13690009", -- 1437c
		x"0009266e", -- 14380
		x"fff8377c", -- 14384
		x"0001002c", -- 14388
		x"4a2a000f", -- 1438c
		x"67000010", -- 14390
		x"286e0008", -- 14394
		x"28bc0000", -- 14398
		x"00016000", -- 1439c
		x"00b22f2e", -- 143a0
		x"000c2f2e", -- 143a4
		x"00084eb9", -- 143a8
		x"00011f7c", -- 143ac
		x"206e0008", -- 143b0
		x"7005b090", -- 143b4
		x"66000080", -- 143b8
		x"2f2e000c", -- 143bc
		x"2f2e0008", -- 143c0
		x"4ebaf6c0", -- 143c4
		x"206e0008", -- 143c8
		x"7010b090", -- 143cc
		x"57c06700", -- 143d0
		x"0014206e", -- 143d4
		x"0008700c", -- 143d8
		x"b09057c0", -- 143dc
		x"67000006", -- 143e0
		x"60000038", -- 143e4
		x"2f2e000c", -- 143e8
		x"2f2e0008", -- 143ec
		x"4ebafe18", -- 143f0
		x"206effe4", -- 143f4
		x"7002b050", -- 143f8
		x"6600000c", -- 143fc
		x"1d680003", -- 14400
		x"fffd6000", -- 14404
		x"00081d7c", -- 14408
		x"0000fffd", -- 1440c
		x"206effe8", -- 14410
		x"116efffd", -- 14414
		x"00076000", -- 14418
		x"001a206e", -- 1441c
		x"000820bc", -- 14420
		x"00000001", -- 14424
		x"2f2e000c", -- 14428
		x"3f3c000d", -- 1442c
		x"4eb90001", -- 14430
		x"18806000", -- 14434
		x"001a206e", -- 14438
		x"000820bc", -- 1443c
		x"00000001", -- 14440
		x"2f2e000c", -- 14444
		x"3f3c0008", -- 14448
		x"4eb90001", -- 1444c
		x"18804e5e", -- 14450
		x"205f504f", -- 14454
		x"4ed00000", -- 14458
		x"4e56fff8", -- 1445c
		x"2d6e000c", -- 14460
		x"fffc206e", -- 14464
		x"fffc2268", -- 14468
		x"00482d69", -- 1446c
		x"0044fff8", -- 14470
		x"7001b068", -- 14474
		x"002c6600", -- 14478
		x"0020226e", -- 1447c
		x"fff80829", -- 14480
		x"0007000d", -- 14484
		x"56c04400", -- 14488
		x"4a006700", -- 1448c
		x"000c206e", -- 14490
		x"00084290", -- 14494
		x"6000002e", -- 14498
		x"206efff8", -- 1449c
		x"08280003", -- 144a0
		x"000b56c0", -- 144a4
		x"44004a00", -- 144a8
		x"67000010", -- 144ac
		x"226e0008", -- 144b0
		x"22bc0000", -- 144b4
		x"00046000", -- 144b8
		x"000c206e", -- 144bc
		x"000820bc", -- 144c0
		x"00000003", -- 144c4
		x"4e5e205f", -- 144c8
		x"504f4ed0", -- 144cc
		x"00004e56", -- 144d0
		x"fffe3d7c", -- 144d4
		x"0006fffe", -- 144d8
		x"558f2f2e", -- 144dc
		x"000c486e", -- 144e0
		x"fffe3f3c", -- 144e4
		x"00064227", -- 144e8
		x"42274eb9", -- 144ec
		x"00012454", -- 144f0
		x"4a1f6700", -- 144f4
		x"000c206e", -- 144f8
		x"00084290", -- 144fc
		x"6000001a", -- 14500
		x"206e0008", -- 14504
		x"20bc0000", -- 14508
		x"00012f2e", -- 1450c
		x"000c3f3c", -- 14510
		x"00084eb9", -- 14514
		x"00011880", -- 14518
		x"4e5e205f", -- 1451c
		x"504f4ed0", -- 14520
		x"4e750000", -- 14524
		x"4e56ffec", -- 14528
		x"598f3f2e", -- 1452c
		x"00084eb9", -- 14530
		x"00011a02", -- 14534
		x"2d5ffff8", -- 14538
		x"2d6efff8", -- 1453c
		x"fff0206e", -- 14540
		x"fff04a28", -- 14544
		x"004c6700", -- 14548
		x"002c2f28", -- 1454c
		x"004e1f28", -- 14550
		x"004d4eb9", -- 14554
		x"00011d94", -- 14558
		x"3f2e0008", -- 1455c
		x"4eb90001", -- 14560
		x"1f28206e", -- 14564
		x"fff04228", -- 14568
		x"004c2268", -- 1456c
		x"0040137c", -- 14570
		x"00010007", -- 14574
		x"2d7cffff", -- 14578
		x"fffffff4", -- 1457c
		x"52aefff4", -- 14580
		x"206efff0", -- 14584
		x"202efff4", -- 14588
		x"e5804ab0", -- 1458c
		x"08006700", -- 14590
		x"004e202e", -- 14594
		x"fff4e580", -- 14598
		x"2d700800", -- 1459c
		x"fffc202e", -- 145a0
		x"fff4e580", -- 145a4
		x"42b00800", -- 145a8
		x"2d6efffc", -- 145ac
		x"ffec2f2e", -- 145b0
		x"fffc3f3c", -- 145b4
		x"000c4eb9", -- 145b8
		x"00011880", -- 145bc
		x"206effec", -- 145c0
		x"317c0003", -- 145c4
		x"002c4a28", -- 145c8
		x"004c6700", -- 145cc
		x"00124aa8", -- 145d0
		x"00286704", -- 145d4
		x"2f280028", -- 145d8
		x"22680024", -- 145dc
		x"4e910cae", -- 145e0
		x"00000007", -- 145e4
		x"fff46d94", -- 145e8
		x"4e5e205f", -- 145ec
		x"544f4ed0", -- 145f0
		x"00004e56", -- 145f4
		x"0000598f", -- 145f8
		x"3f2e0008", -- 145fc
		x"4eb90001", -- 14600
		x"1a02205f", -- 14604
		x"20680044", -- 14608
		x"08280003", -- 1460c
		x"000b56c0", -- 14610
		x"44004a00", -- 14614
		x"6700000c", -- 14618
		x"3f2e0008", -- 1461c
		x"4eb90001", -- 14620
		x"236a3f2e", -- 14624
		x"00084eb9", -- 14628
		x"0001227e", -- 1462c
		x"3f2e0008", -- 14630
		x"4ebafef2", -- 14634
		x"4e5e205f", -- 14638
		x"544f4ed0", -- 1463c
		x"00004e56", -- 14640
		x"ffec2d6e", -- 14644
		x"000cfff4", -- 14648
		x"206e000c", -- 1464c
		x"41e80044", -- 14650
		x"2d48fff0", -- 14654
		x"206efff4", -- 14658
		x"42680030", -- 1465c
		x"4268002e", -- 14660
		x"4268002c", -- 14664
		x"226efff0", -- 14668
		x"4229000e", -- 1466c
		x"42690012", -- 14670
		x"4ca81e00", -- 14674
		x"002448ae", -- 14678
		x"1e00fff8", -- 1467c
		x"4aaefff8", -- 14680
		x"56c0226e", -- 14684
		x"fff00200", -- 14688
		x"ff011340", -- 1468c
		x"0008237c", -- 14690
		x"000145f6", -- 14694
		x"003242a9", -- 14698
		x"0036598f", -- 1469c
		x"3f104eb9", -- 146a0
		x"00011a02", -- 146a4
		x"206efff0", -- 146a8
		x"215f0004", -- 146ac
		x"4aa80004", -- 146b0
		x"66000028", -- 146b4
		x"2f2e000c", -- 146b8
		x"3f3c0005", -- 146bc
		x"4eb90001", -- 146c0
		x"1880206e", -- 146c4
		x"fff4317c", -- 146c8
		x"0003002c", -- 146cc
		x"226e0008", -- 146d0
		x"22bc0000", -- 146d4
		x"00016000", -- 146d8
		x"0066206e", -- 146dc
		x"fff02d68", -- 146e0
		x"0004ffec", -- 146e4
		x"226effec", -- 146e8
		x"246efff4", -- 146ec
		x"302a0002", -- 146f0
		x"48c0e580", -- 146f4
		x"4ab10800", -- 146f8
		x"67000028", -- 146fc
		x"2f2e000c", -- 14700
		x"3f3c0001", -- 14704
		x"4eb90001", -- 14708
		x"1880206e", -- 1470c
		x"fff4317c", -- 14710
		x"0003002c", -- 14714
		x"226e0008", -- 14718
		x"22bc0000", -- 1471c
		x"00016000", -- 14720
		x"001e206e", -- 14724
		x"ffec226e", -- 14728
		x"fff43029", -- 1472c
		x"000248c0", -- 14730
		x"e58021ae", -- 14734
		x"000c0800", -- 14738
		x"246e0008", -- 1473c
		x"42924e5e", -- 14740
		x"205f504f", -- 14744
		x"4ed00000", -- 14748
		x"4e56fff4", -- 1474c
		x"2f2e0008", -- 14750
		x"486efffc", -- 14754
		x"4ebafee8", -- 14758
		x"4aaefffc", -- 1475c
		x"6600000c", -- 14760
		x"2f2e0008", -- 14764
		x"4eb90001", -- 14768
		x"2e7c2d6e", -- 1476c
		x"0008fff4", -- 14770
		x"206efff4", -- 14774
		x"4a280052", -- 14778
		x"67000046", -- 1477c
		x"598f3f10", -- 14780
		x"4eb90001", -- 14784
		x"1a022d5f", -- 14788
		x"fff8206e", -- 1478c
		x"fff82068", -- 14790
		x"00400828", -- 14794
		x"00060003", -- 14798
		x"56c04400", -- 1479c
		x"4a006600", -- 147a0
		x"000460e6", -- 147a4
		x"206efff4", -- 147a8
		x"3f10226e", -- 147ac
		x"fff84aa9", -- 147b0
		x"00566704", -- 147b4
		x"2f290056", -- 147b8
		x"22690052", -- 147bc
		x"4e9160b0", -- 147c0
		x"4e5e2e9f", -- 147c4
		x"4e750000", -- 147c8
		x"4e56fffa", -- 147cc
		x"558f2f2e", -- 147d0
		x"000c486e", -- 147d4
		x"fffe3f3c", -- 147d8
		x"00034227", -- 147dc
		x"42274eb9", -- 147e0
		x"00012454", -- 147e4
		x"4a1f6700", -- 147e8
		x"0022206e", -- 147ec
		x"00084290", -- 147f0
		x"2d6e000c", -- 147f4
		x"fffa206e", -- 147f8
		x"fffa316e", -- 147fc
		x"fffe002e", -- 14800
		x"2168006c", -- 14804
		x"00326000", -- 14808
		x"001a206e", -- 1480c
		x"000820bc", -- 14810
		x"00000001", -- 14814
		x"2f2e000c", -- 14818
		x"3f3c0008", -- 1481c
		x"4eb90001", -- 14820
		x"18804e5e", -- 14824
		x"205f504f", -- 14828
		x"4ed00000", -- 1482c
		x"4e560000", -- 14830
		x"206e0008", -- 14834
		x"20bc0000", -- 14838
		x"00014e5e", -- 1483c
		x"205f504f", -- 14840
		x"4ed00000", -- 14844
		x"4e56fff4", -- 14848
		x"206e0008", -- 1484c
		x"42902d6e", -- 14850
		x"000cfffc", -- 14854
		x"206efffc", -- 14858
		x"43e80044", -- 1485c
		x"2d49fff8", -- 14860
		x"226efff8", -- 14864
		x"2d690004", -- 14868
		x"fff4317c", -- 1486c
		x"0003002c", -- 14870
		x"4a290008", -- 14874
		x"67000012", -- 14878
		x"4aa80028", -- 1487c
		x"67042f28", -- 14880
		x"00282468", -- 14884
		x"00244e92", -- 14888
		x"206efff4", -- 1488c
		x"226efffc", -- 14890
		x"30290002", -- 14894
		x"48c0e580", -- 14898
		x"42b00800", -- 1489c
		x"4e5e205f", -- 148a0
		x"504f4ed0", -- 148a4
		x"00004e56", -- 148a8
		x"00002f2e", -- 148ac
		x"000c3f3c", -- 148b0
		x"00034eb9", -- 148b4
		x"00011880", -- 148b8
		x"206e0008", -- 148bc
		x"42904e5e", -- 148c0
		x"205f504f", -- 148c4
		x"4ed00000", -- 148c8
		x"4e560000", -- 148cc
		x"2f2e000c", -- 148d0
		x"3f3c000b", -- 148d4
		x"4eb90001", -- 148d8
		x"1880206e", -- 148dc
		x"00084290", -- 148e0
		x"4e5e205f", -- 148e4
		x"504f4ed0", -- 148e8
		x"00004e56", -- 148ec
		x"0000206e", -- 148f0
		x"000c3f10", -- 148f4
		x"4ebafc2e", -- 148f8
		x"206e0008", -- 148fc
		x"42904e5e", -- 14900
		x"205f504f", -- 14904
		x"4ed04e75", -- 14908
		x"00004e56", -- 1490c
		x"ffd42f2d", -- 14910
		x"fff62f0e", -- 14914
		x"487a01dc", -- 14918
		x"2b4ffff6", -- 1491c
		x"42aeffe4", -- 14920
		x"598f3f2e", -- 14924
		x"00084eb9", -- 14928
		x"00011a02", -- 1492c
		x"2d5ffffc", -- 14930
		x"2d6efffc", -- 14934
		x"ffe0206e", -- 14938
		x"ffe02d68", -- 1493c
		x"0044ffdc", -- 14940
		x"422effef", -- 14944
		x"42aefff0", -- 14948
		x"206effe0", -- 1494c
		x"202efff0", -- 14950
		x"e5802d70", -- 14954
		x"0800fff8", -- 14958
		x"4aaefff8", -- 1495c
		x"6700003e", -- 14960
		x"2d6efff8", -- 14964
		x"ffd8226e", -- 14968
		x"ffd845e9", -- 1496c
		x"00442d4a", -- 14970
		x"ffd47001", -- 14974
		x"b069002c", -- 14978
		x"66000022", -- 1497c
		x"246effd4", -- 14980
		x"4a2a000e", -- 14984
		x"67000016", -- 14988
		x"1d7c0001", -- 1498c
		x"ffef206e", -- 14990
		x"ffd43028", -- 14994
		x"001048c0", -- 14998
		x"2d40ffe4", -- 1499c
		x"52aefff0", -- 149a0
		x"102effef", -- 149a4
		x"66000010", -- 149a8
		x"7007b0ae", -- 149ac
		x"fff05dc0", -- 149b0
		x"6d000004", -- 149b4
		x"60924a2e", -- 149b8
		x"ffef6600", -- 149bc
		x"00b0206e", -- 149c0
		x"ffdc7040", -- 149c4
		x"b0280009", -- 149c8
		x"660000a2", -- 149cc
		x"206effdc", -- 149d0
		x"70001028", -- 149d4
		x"00177200", -- 149d8
		x"12280001", -- 149dc
		x"904148c0", -- 149e0
		x"2d40fff0", -- 149e4
		x"42aefff4", -- 149e8
		x"7001b0ae", -- 149ec
		x"fff06700", -- 149f0
		x"00287007", -- 149f4
		x"b0aefff4", -- 149f8
		x"6f00001e", -- 149fc
		x"598f2f2e", -- 14a00
		x"fff02f3c", -- 14a04
		x"00000001", -- 14a08
		x"4eb90001", -- 14a0c
		x"4b662d5f", -- 14a10
		x"fff052ae", -- 14a14
		x"fff460d0", -- 14a18
		x"206effe0", -- 14a1c
		x"202efff4", -- 14a20
		x"e5802d70", -- 14a24
		x"0800fff8", -- 14a28
		x"4aaefff8", -- 14a2c
		x"6700003e", -- 14a30
		x"2d6efff8", -- 14a34
		x"ffd8226e", -- 14a38
		x"ffd845e9", -- 14a3c
		x"00442d4a", -- 14a40
		x"ffd47002", -- 14a44
		x"b069002c", -- 14a48
		x"66000022", -- 14a4c
		x"246effd4", -- 14a50
		x"4a2a000e", -- 14a54
		x"67000016", -- 14a58
		x"1d7c0001", -- 14a5c
		x"ffef206e", -- 14a60
		x"ffd43028", -- 14a64
		x"001048c0", -- 14a68
		x"2d40ffe4", -- 14a6c
		x"4a2effef", -- 14a70
		x"6700003a", -- 14a74
		x"4aaeffe4", -- 14a78
		x"67000032", -- 14a7c
		x"598f206e", -- 14a80
		x"ffdc7000", -- 14a84
		x"10280009", -- 14a88
		x"2f002f2e", -- 14a8c
		x"ffe44eb9", -- 14a90
		x"00014b46", -- 14a94
		x"201fb0ae", -- 14a98
		x"ffe46600", -- 14a9c
		x"00102f2e", -- 14aa0
		x"fff84eb9", -- 14aa4
		x"00012e7c", -- 14aa8
		x"6000003a", -- 14aac
		x"4a2effef", -- 14ab0
		x"67000028", -- 14ab4
		x"2f2efff8", -- 14ab8
		x"3f3c0004", -- 14abc
		x"4eb90001", -- 14ac0
		x"1880206e", -- 14ac4
		x"fff8117c", -- 14ac8
		x"ff010053", -- 14acc
		x"2f2efff8", -- 14ad0
		x"4eb90001", -- 14ad4
		x"2e7c6000", -- 14ad8
		x"000c3f2e", -- 14adc
		x"00084eb9", -- 14ae0
		x"000145f6", -- 14ae4
		x"2b6f0008", -- 14ae8
		x"fff6defc", -- 14aec
		x"000c4efa", -- 14af0
		x"00122c5f", -- 14af4
		x"2b5ffff6", -- 14af8
		x"3f2e0008", -- 14afc
		x"4eb90001", -- 14b00
		x"45f64e5e", -- 14b04
		x"205f544f", -- 14b08
		x"4ed04e75", -- 14b0c
		x"4ef90000", -- 14b10
		x"526e205f", -- 14b14
		x"2278fed4", -- 14b18
		x"22690010", -- 14b1c
		x"235f0012", -- 14b20
		x"48690012", -- 14b24
		x"2f084ef9", -- 14b28
		x"0000521e", -- 14b2c
		x"205f2278", -- 14b30
		x"fed42269", -- 14b34
		x"00104869", -- 14b38
		x"00122f08", -- 14b3c
		x"4ef90000", -- 14b40
		x"5258205f", -- 14b44
		x"201f809f", -- 14b48
		x"2e804ed0", -- 14b4c
		x"205f201f", -- 14b50
		x"c09f2e80", -- 14b54
		x"4ed0205f", -- 14b58
		x"201f221f", -- 14b5c
		x"e1a92e81", -- 14b60
		x"4ed0205f", -- 14b64
		x"201f221f", -- 14b68
		x"e0a92e81", -- 14b6c
		x"4ed04e56", -- 14b70
		x"fffc4aae", -- 14b74
		x"00086e0a", -- 14b78
		x"0caef332", -- 14b7c
		x"a9600008", -- 14b80
		x"60222d7c", -- 14b84
		x"00000001", -- 14b88
		x"fffc202e", -- 14b8c
		x"fffcb0ae", -- 14b90
		x"00086c08", -- 14b94
		x"e3802d40", -- 14b98
		x"fffc60ee", -- 14b9c
		x"202efffc", -- 14ba0
		x"b0ae0008", -- 14ba4
		x"57c00200", -- 14ba8
		x"00011d40", -- 14bac
		x"000c4e5e", -- 14bb0
		x"2e9f4e75", -- 14bb4
		x"225f205f", -- 14bb8
		x"4a1f7000", -- 14bbc
		x"10106f10", -- 14bc0
		x"45f00801", -- 14bc4
		x"7220b222", -- 14bc8
		x"66045380", -- 14bcc
		x"6ef81080", -- 14bd0
		x"4ed14e75", -- 14bd4
		x"01360002", -- 14bd8
		x"03010004", -- 14bdc
		x"00160003", -- 14be0
		x"002a0001", -- 14be4
		x"00520001", -- 14be8
		x"1f7c0002", -- 14bec
		x"03010002", -- 14bf0
		x"00660003", -- 14bf4
		x"002a0001", -- 14bf8
		x"00520001", -- 14bfc
		x"2ff60102", -- 14c00
		x"08010007", -- 14c04
		x"006a0001", -- 14c08
		x"00520004", -- 14c0c
		x"00160003", -- 14c10
		x"00920005", -- 14c14
		x"00920006", -- 14c18
		x"00920008", -- 14c1c
		x"00920009", -- 14c20
		x"009e0001", -- 14c24
		x"4d3a0103", -- 14c28
		x"03010003", -- 14c2c
		x"01420004", -- 14c30
		x"01420000", -- 14c34
		x"014e0001", -- 14c38
		x"4f4c0300", -- 14c3c
		x"00160102", -- 14c40
		x"08010008", -- 14c44
		x"00ca0009", -- 14c48
		x"009e0001", -- 14c4c
		x"00520004", -- 14c50
		x"00920007", -- 14c54
		x"00920003", -- 14c58
		x"00920005", -- 14c5c
		x"00920006", -- 14c60
		x"00920001", -- 14c64
		x"4ddc0003", -- 14c68
		x"01010000", -- 14c6c
		x"00520001", -- 14c70
		x"48cc0002", -- 14c74
		x"08020005", -- 14c78
		x"00f20001", -- 14c7c
		x"00520008", -- 14c80
		x"00920009", -- 14c84
		x"00920004", -- 14c88
		x"00920007", -- 14c8c
		x"00920003", -- 14c90
		x"00920006", -- 14c94
		x"00920001", -- 14c98
		x"47cc0001", -- 14c9c
		x"1f7c0102", -- 14ca0
		x"08010008", -- 14ca4
		x"00ca0009", -- 14ca8
		x"009e0001", -- 14cac
		x"00520004", -- 14cb0
		x"00920007", -- 14cb4
		x"00920003", -- 14cb8
		x"00920005", -- 14cbc
		x"00920006", -- 14cc0
		x"00920001", -- 14cc4
		x"4ddc0102", -- 14cc8
		x"08010003", -- 14ccc
		x"011a0007", -- 14cd0
		x"01260001", -- 14cd4
		x"00520005", -- 14cd8
		x"00920008", -- 14cdc
		x"00920009", -- 14ce0
		x"00920004", -- 14ce4
		x"00920006", -- 14ce8
		x"00920001", -- 14cec
		x"4efe0003", -- 14cf0
		x"01010000", -- 14cf4
		x"01320001", -- 14cf8
		x"48480003", -- 14cfc
		x"01010000", -- 14d00
		x"006a0001", -- 14d04
		x"48300200", -- 14d08
		x"00000003", -- 14d0c
		x"01010000", -- 14d10
		x"00520001", -- 14d14
		x"48aa0003", -- 14d18
		x"01010000", -- 14d1c
		x"01320001", -- 14d20
		x"48480003", -- 14d24
		x"01030000", -- 14d28
		x"01320001", -- 14d2c
		x"205a0001", -- 14d30
		x"203a0001", -- 14d34
		x"48ee0096", -- 14d38
		x"00030302", -- 14d3c
		x"0002001a", -- 14d40
		x"0006001e", -- 14d44
		x"0000003a", -- 14d48
		x"0001309c", -- 14d4c
		x"00011f7c", -- 14d50
		x"03000002", -- 14d54
		x"00030402", -- 14d58
		x"0013003e", -- 14d5c
		x"00050052", -- 14d60
		x"0001003a", -- 14d64
		x"0000003a", -- 14d68
		x"00013360", -- 14d6c
		x"00011f7c", -- 14d70
		x"02000000", -- 14d74
		x"00030202", -- 14d78
		x"0001003a", -- 14d7c
		x"0000003a", -- 14d80
		x"00013460", -- 14d84
		x"00011f7c", -- 14d88
		x"00030301", -- 14d8c
		x"000a0066", -- 14d90
		x"0001003a", -- 14d94
		x"0000007a", -- 14d98
		x"00013a86", -- 14d9c
		x"00030202", -- 14da0
		x"0001003a", -- 14da4
		x"0000003a", -- 14da8
		x"000137f0", -- 14dac
		x"00011f7c", -- 14db0
		x"00030402", -- 14db4
		x"00050052", -- 14db8
		x"0006003e", -- 14dbc
		x"0001003a", -- 14dc0
		x"0000003a", -- 14dc4
		x"00013c50", -- 14dc8
		x"00011f7c", -- 14dcc
		x"00030101", -- 14dd0
		x"0000003a", -- 14dd4
		x"000148aa", -- 14dd8
		x"01160003", -- 14ddc
		x"01010000", -- 14de0
		x"000e0001", -- 14de4
		x"3cbe0003", -- 14de8
		x"04020002", -- 14dec
		x"002a0005", -- 14df0
		x"002e0006", -- 14df4
		x"004e0000", -- 14df8
		x"00660001", -- 14dfc
		x"3df80001", -- 14e00
		x"1f7c0300", -- 14e04
		x"000e0003", -- 14e08
		x"0601000b", -- 14e0c
		x"006a000c", -- 14e10
		x"007e000d", -- 14e14
		x"0092000a", -- 14e18
		x"00aa0001", -- 14e1c
		x"00660000", -- 14e20
		x"00be0001", -- 14e24
		x"3a860003", -- 14e28
		x"03020005", -- 14e2c
		x"002e0001", -- 14e30
		x"00660000", -- 14e34
		x"00660001", -- 14e38
		x"3fb80001", -- 14e3c
		x"1f7c0200", -- 14e40
		x"00000003", -- 14e44
		x"02020005", -- 14e48
		x"002e0000", -- 14e4c
		x"00d60001", -- 14e50
		x"40460001", -- 14e54
		x"1f7c0003", -- 14e58
		x"02020005", -- 14e5c
		x"002e0000", -- 14e60
		x"00d60001", -- 14e64
		x"420a0001", -- 14e68
		x"1f7c0002", -- 14e6c
		x"03020002", -- 14e70
		x"00e60003", -- 14e74
		x"00ea0001", -- 14e78
		x"00660001", -- 14e7c
		x"41ec0001", -- 14e80
		x"2ff60003", -- 14e84
		x"02020001", -- 14e88
		x"00660000", -- 14e8c
		x"00d60001", -- 14e90
		x"37f00001", -- 14e94
		x"1f7c0003", -- 14e98
		x"03020005", -- 14e9c
		x"002e0001", -- 14ea0
		x"00660000", -- 14ea4
		x"00d60001", -- 14ea8
		x"3c500001", -- 14eac
		x"1f7c0003", -- 14eb0
		x"02010014", -- 14eb4
		x"010a0000", -- 14eb8
		x"00660001", -- 14ebc
		x"423a0300", -- 14ec0
		x"00920003", -- 14ec4
		x"04020002", -- 14ec8
		x"01060005", -- 14ecc
		x"002e0001", -- 14ed0
		x"00660000", -- 14ed4
		x"00d60001", -- 14ed8
		x"42e40001", -- 14edc
		x"1f7c0300", -- 14ee0
		x"00ea0003", -- 14ee4
		x"01010000", -- 14ee8
		x"000e0001", -- 14eec
		x"3de40003", -- 14ef0
		x"01010000", -- 14ef4
		x"00660001", -- 14ef8
		x"48aa0042", -- 14efc
		x"00030501", -- 14f00
		x"000e001e", -- 14f04
		x"0011001e", -- 14f08
		x"0012001e", -- 14f0c
		x"0001002a", -- 14f10
		x"0000002e", -- 14f14
		x"00013a86", -- 14f18
		x"00030101", -- 14f1c
		x"0000002a", -- 14f20
		x"00011f7c", -- 14f24
		x"02000000", -- 14f28
		x"00030202", -- 14f2c
		x"00050002", -- 14f30
		x"0000002a", -- 14f34
		x"00013c50", -- 14f38
		x"00011f7c", -- 14f3c
		x"00030101", -- 14f40
		x"0000002a", -- 14f44
		x"000148aa", -- 14f48
		x"003a0003", -- 14f4c
		x"02010000", -- 14f50
		x"00120000", -- 14f54
		x"00220001", -- 14f58
		x"445c0002", -- 14f5c
		x"02010006", -- 14f60
		x"00260001", -- 14f64
		x"00220001", -- 14f68
		x"207a0200", -- 14f6c
		x"00000003", -- 14f70
		x"02020001", -- 14f74
		x"00220000", -- 14f78
		x"00220001", -- 14f7c
		x"44d20001", -- 14f80
		x"1f7c0003", -- 14f84
		x"01010000", -- 14f88
		x"00220001", -- 14f8c
		x"48aaffff", -- 14f90
		x"c3b3a6b0", -- 14f94
		x"ffff48e7", -- 14f98
		x"fffe2a78", -- 14f9c
		x"fed46100", -- 14fa0
		x"00ec4284", -- 14fa4
		x"42854286", -- 14fa8
		x"428749f9", -- 14fac
		x"00500000", -- 14fb0
		x"3c3c0004", -- 14fb4
		x"383c008f", -- 14fb8
		x"6176662c", -- 14fbc
		x"49f90050", -- 14fc0
		x"00083c3c", -- 14fc4
		x"0004383c", -- 14fc8
		x"00ff6164", -- 14fcc
		x"661a0c2d", -- 14fd0
		x"0003033f", -- 14fd4
		x"6d1249f9", -- 14fd8
		x"00500100", -- 14fdc
		x"61146608", -- 14fe0
		x"49f90050", -- 14fe4
		x"0200610a", -- 14fe8
		x"4a2d0328", -- 14fec
		x"4cdf7fff", -- 14ff0
		x"4e753c3c", -- 14ff4
		x"0000383c", -- 14ff8
		x"ffff6134", -- 14ffc
		x"662e3c3c", -- 15000
		x"0002383c", -- 15004
		x"ffff6128", -- 15008
		x"66223c3c", -- 1500c
		x"0004383c", -- 15010
		x"ffff611c", -- 15014
		x"66163c3c", -- 15018
		x"0006383c", -- 1501c
		x"ffff6110", -- 15020
		x"660a3c3c", -- 15024
		x"0008383c", -- 15028
		x"06ff6104", -- 1502c
		x"615e4e75", -- 15030
		x"610c56ed", -- 15034
		x"03286154", -- 15038
		x"4a2d0328", -- 1503c
		x"4e7548e7", -- 15040
		x"f4844205", -- 15044
		x"303c8000", -- 15048
		x"32003401", -- 1504c
		x"c2444642", -- 15050
		x"c4443982", -- 15054
		x"60004e71", -- 15058
		x"36346000", -- 1505c
		x"c644b642", -- 15060
		x"661a3401", -- 15064
		x"39826000", -- 15068
		x"4e713634", -- 1506c
		x"6000c644", -- 15070
		x"b6426608", -- 15074
		x"4a40670c", -- 15078
		x"e24860cc", -- 1507c
		x"50c53806", -- 15080
		x"3c023e03", -- 15084
		x"4a054cdf", -- 15088
		x"212f4e75", -- 1508c
		x"4a790050", -- 15090
		x"00004a79", -- 15094
		x"00500008", -- 15098
		x"4e7548e7", -- 1509c
		x"fffe2a78", -- 150a0
		x"fdce2b4f", -- 150a4
		x"00044dfa", -- 150a8
		x"03a841ed", -- 150ac
		x"00142008", -- 150b0
		x"c0bc0000", -- 150b4
		x"00036706", -- 150b8
		x"72049280", -- 150bc
		x"d1c12b48", -- 150c0
		x"000841e8", -- 150c4
		x"00402b48", -- 150c8
		x"000c41e8", -- 150cc
		x"00402b48", -- 150d0
		x"0010422d", -- 150d4
		x"0001422d", -- 150d8
		x"000208ea", -- 150dc
		x"00020003", -- 150e0
		x"082a0002", -- 150e4
		x"00036704", -- 150e8
		x"522d0002", -- 150ec
		x"4a2d0002", -- 150f0
		x"67000348", -- 150f4
		x"610002f6", -- 150f8
		x"66000340", -- 150fc
		x"610005bc", -- 15100
		x"66000338", -- 15104
		x"42844285", -- 15108
		x"42864287", -- 1510c
		x"383c008f", -- 15110
		x"3c3c0002", -- 15114
		x"61000630", -- 15118
		x"66000320", -- 1511c
		x"383c00ff", -- 15120
		x"3c3c0012", -- 15124
		x"61000620", -- 15128
		x"66000310", -- 1512c
		x"383c00c0", -- 15130
		x"3c3c0016", -- 15134
		x"61000610", -- 15138
		x"66000300", -- 1513c
		x"383c00fe", -- 15140
		x"3c3c0018", -- 15144
		x"61000600", -- 15148
		x"660002f0", -- 1514c
		x"383c00ff", -- 15150
		x"3c3c001a", -- 15154
		x"610005f0", -- 15158
		x"660002e0", -- 1515c
		x"383c00ff", -- 15160
		x"3c3c001c", -- 15164
		x"610005e0", -- 15168
		x"660002d0", -- 1516c
		x"383c00ff", -- 15170
		x"3c3c001e", -- 15174
		x"610005d0", -- 15178
		x"660002c0", -- 1517c
		x"4a2d0001", -- 15180
		x"660002b8", -- 15184
		x"42526100", -- 15188
		x"05266100", -- 1518c
		x"052e6100", -- 15190
		x"057a002a", -- 15194
		x"00800019", -- 15198
		x"3e3c001e", -- 1519c
		x"103c0055", -- 151a0
		x"6100049c", -- 151a4
		x"4a2d0001", -- 151a8
		x"66264600", -- 151ac
		x"61000490", -- 151b0
		x"4a2d0001", -- 151b4
		x"661a303c", -- 151b8
		x"01006100", -- 151bc
		x"04824a2d", -- 151c0
		x"0001660c", -- 151c4
		x"46006100", -- 151c8
		x"04764a2d", -- 151cc
		x"00016704", -- 151d0
		x"60000268", -- 151d4
		x"4600e258", -- 151d8
		x"6ce0022a", -- 151dc
		x"003f0017", -- 151e0
		x"002a0080", -- 151e4
		x"0017157c", -- 151e8
		x"00000013", -- 151ec
		x"4201102a", -- 151f0
		x"00116600", -- 151f4
		x"0136157c", -- 151f8
		x"00a50015", -- 151fc
		x"2f3c0000", -- 15200
		x"00044eb9", -- 15204
		x"0000526e", -- 15208
		x"102a0011", -- 1520c
		x"6600011c", -- 15210
		x"102a0015", -- 15214
		x"2f3c0000", -- 15218
		x"00044eb9", -- 1521c
		x"0000526e", -- 15220
		x"123c008a", -- 15224
		x"022a003f", -- 15228
		x"0017002a", -- 1522c
		x"00400017", -- 15230
		x"157c00ff", -- 15234
		x"0013102a", -- 15238
		x"0011b001", -- 1523c
		x"660000ec", -- 15240
		x"123c008e", -- 15244
		x"15400015", -- 15248
		x"2f3c0000", -- 1524c
		x"00044eb9", -- 15250
		x"0000526e", -- 15254
		x"102a0011", -- 15258
		x"b0016600", -- 1525c
		x"00ce123c", -- 15260
		x"008e343c", -- 15264
		x"00061540", -- 15268
		x"00152f3c", -- 1526c
		x"00000004", -- 15270
		x"4eb90000", -- 15274
		x"526e102a", -- 15278
		x"0011b001", -- 1527c
		x"660000ac", -- 15280
		x"51caffe4", -- 15284
		x"123c008c", -- 15288
		x"343c0006", -- 1528c
		x"15400015", -- 15290
		x"2f3c0000", -- 15294
		x"00044eb9", -- 15298
		x"0000526e", -- 1529c
		x"102a0011", -- 152a0
		x"b0016600", -- 152a4
		x"008651ca", -- 152a8
		x"ffe4123c", -- 152ac
		x"00841540", -- 152b0
		x"00152f3c", -- 152b4
		x"00000004", -- 152b8
		x"4eb90000", -- 152bc
		x"526e102a", -- 152c0
		x"0011b001", -- 152c4
		x"66000064", -- 152c8
		x"123c00c4", -- 152cc
		x"15400015", -- 152d0
		x"2f3c0000", -- 152d4
		x"00044eb9", -- 152d8
		x"0000526e", -- 152dc
		x"102a0011", -- 152e0
		x"b0016600", -- 152e4
		x"0046123c", -- 152e8
		x"00ca343c", -- 152ec
		x"000f102a", -- 152f0
		x"00152f3c", -- 152f4
		x"00000004", -- 152f8
		x"4eb90000", -- 152fc
		x"526e51ca", -- 15300
		x"ffee102a", -- 15304
		x"0011b001", -- 15308
		x"6620157c", -- 1530c
		x"00ff0011", -- 15310
		x"123c000a", -- 15314
		x"2f3c0000", -- 15318
		x"00044eb9", -- 1531c
		x"0000526e", -- 15320
		x"102a0011", -- 15324
		x"b0016602", -- 15328
		x"600850ed", -- 1532c
		x"00016000", -- 15330
		x"010a157c", -- 15334
		x"00010001", -- 15338
		x"2878fed4", -- 1533c
		x"4a2c033f", -- 15340
		x"670000f8", -- 15344
		x"266d0010", -- 15348
		x"61000364", -- 1534c
		x"610a6100", -- 15350
		x"03526104", -- 15354
		x"60000092", -- 15358
		x"615c6112", -- 1535c
		x"6162610e", -- 15360
		x"6168610a", -- 15364
		x"616e6106", -- 15368
		x"61746102", -- 1536c
		x"4e756100", -- 15370
		x"00ee6102", -- 15374
		x"4e754a2d", -- 15378
		x"00016702", -- 1537c
		x"6136206d", -- 15380
		x"0008226d", -- 15384
		x"000c4242", -- 15388
		x"b3886702", -- 1538c
		x"61205842", -- 15390
		x"4a2d0000", -- 15394
		x"67080c42", -- 15398
		x"002066ec", -- 1539c
		x"60060c42", -- 153a0
		x"004066e4", -- 153a4
		x"4a2d0001", -- 153a8
		x"66000090", -- 153ac
		x"4e7550ed", -- 153b0
		x"00014e75", -- 153b4
		x"4e75203c", -- 153b8
		x"12345678", -- 153bc
		x"6000025c", -- 153c0
		x"203cf0f0", -- 153c4
		x"f0f06000", -- 153c8
		x"0252203c", -- 153cc
		x"ff00ff00", -- 153d0
		x"60000248", -- 153d4
		x"203caaaa", -- 153d8
		x"aaab6000", -- 153dc
		x"023e203c", -- 153e0
		x"5a5a5a59", -- 153e4
		x"60000234", -- 153e8
		x"6102604e", -- 153ec
		x"610002cc", -- 153f0
		x"6642157c", -- 153f4
		x"00000017", -- 153f8
		x"157c0090", -- 153fc
		x"00192f3c", -- 15400
		x"00000064", -- 15404
		x"4eb90000", -- 15408
		x"526e157c", -- 1540c
		x"00800019", -- 15410
		x"157c0040", -- 15414
		x"0017157c", -- 15418
		x"005e0015", -- 1541c
		x"157c0040", -- 15420
		x"0017157c", -- 15424
		x"00980015", -- 15428
		x"157c00c0", -- 1542c
		x"0017157c", -- 15430
		x"00000015", -- 15434
		x"4a2d0001", -- 15438
		x"4e752a78", -- 1543c
		x"fdce2e6d", -- 15440
		x"00046100", -- 15444
		x"02764a2d", -- 15448
		x"00014cdf", -- 1544c
		x"7fff4e75", -- 15450
		x"2a78fdce", -- 15454
		x"50ed0001", -- 15458
		x"2e6d0004", -- 1545c
		x"60e86100", -- 15460
		x"025a6100", -- 15464
		x"02c048e7", -- 15468
		x"fff0206d", -- 1546c
		x"0008323c", -- 15470
		x"000c203c", -- 15474
		x"0000000f", -- 15478
		x"61000170", -- 1547c
		x"4a2d0000", -- 15480
		x"670c323c", -- 15484
		x"0008d1fc", -- 15488
		x"00000040", -- 1548c
		x"6006d1fc", -- 15490
		x"00000010", -- 15494
		x"61000160", -- 15498
		x"157c0000", -- 1549c
		x"0017157c", -- 154a0
		x"00ff0013", -- 154a4
		x"157c0082", -- 154a8
		x"0019226d", -- 154ac
		x"000c103c", -- 154b0
		x"00094a2d", -- 154b4
		x"00006704", -- 154b8
		x"103c000d", -- 154bc
		x"15400003", -- 154c0
		x"2f3c0000", -- 154c4
		x"00324eb9", -- 154c8
		x"0000526e", -- 154cc
		x"157c0000", -- 154d0
		x"00034a2d", -- 154d4
		x"0000670c", -- 154d8
		x"103c0006", -- 154dc
		x"157c0080", -- 154e0
		x"00196008", -- 154e4
		x"610000d4", -- 154e8
		x"103c000a", -- 154ec
		x"15400003", -- 154f0
		x"2f3c0000", -- 154f4
		x"00324eb9", -- 154f8
		x"0000526e", -- 154fc
		x"157c0000", -- 15500
		x"00034a2d", -- 15504
		x"00006612", -- 15508
		x"610000b0", -- 1550c
		x"d1fc0000", -- 15510
		x"00102008", -- 15514
		x"20492240", -- 15518
		x"600691fc", -- 1551c
		x"00000030", -- 15520
		x"323c0008", -- 15524
		x"203c0000", -- 15528
		x"000f6100", -- 1552c
		x"00be4a2d", -- 15530
		x"0000670c", -- 15534
		x"323c000c", -- 15538
		x"d1fc0000", -- 1553c
		x"00406006", -- 15540
		x"d1fc0000", -- 15544
		x"00106100", -- 15548
		x"00ae103c", -- 1554c
		x"00014a2d", -- 15550
		x"0000670c", -- 15554
		x"103c000e", -- 15558
		x"157c0082", -- 1555c
		x"0019600a", -- 15560
		x"61000070", -- 15564
		x"157c0080", -- 15568
		x"00191540", -- 1556c
		x"00032f3c", -- 15570
		x"00000032", -- 15574
		x"4eb90000", -- 15578
		x"526e157c", -- 1557c
		x"00000003", -- 15580
		x"157c0080", -- 15584
		x"0019103c", -- 15588
		x"00054a2d", -- 1558c
		x"00006606", -- 15590
		x"103c0002", -- 15594
		x"613c1540", -- 15598
		x"00032f3c", -- 1559c
		x"00000032", -- 155a0
		x"4eb90000", -- 155a4
		x"526e157c", -- 155a8
		x"00000003", -- 155ac
		x"4a2d0000", -- 155b0
		x"6602611e", -- 155b4
		x"4cdf0fff", -- 155b8
		x"4e75082a", -- 155bc
		x"00020011", -- 155c0
		x"670e12ea", -- 155c4
		x"0015b3cb", -- 155c8
		x"6ff008ed", -- 155cc
		x"00070001", -- 155d0
		x"4e75082a", -- 155d4
		x"00030011", -- 155d8
		x"670e1559", -- 155dc
		x"0015b3cb", -- 155e0
		x"6ff008ed", -- 155e4
		x"00000001", -- 155e8
		x"4e7548e7", -- 155ec
		x"8040227c", -- 155f0
		x"00500000", -- 155f4
		x"600a48e7", -- 155f8
		x"8040227c", -- 155fc
		x"00500008", -- 15600
		x"4a2d0000", -- 15604
		x"6706e248", -- 15608
		x"08c10001", -- 1560c
		x"4a5122c8", -- 15610
		x"32c032c1", -- 15614
		x"4cdf0201", -- 15618
		x"4e7548e7", -- 1561c
		x"80c0206d", -- 15620
		x"0008226d", -- 15624
		x"000c20c0", -- 15628
		x"e298b1c9", -- 1562c
		x"6df84680", -- 15630
		x"e39822c0", -- 15634
		x"b3cb6df8", -- 15638
		x"4cdf0301", -- 1563c
		x"4e7548e7", -- 15640
		x"f0006100", -- 15644
		x"00c6157c", -- 15648
		x"00400017", -- 1564c
		x"12070601", -- 15650
		x"00201541", -- 15654
		x"00150601", -- 15658
		x"00201541", -- 1565c
		x"0015157c", -- 15660
		x"00000017", -- 15664
		x"363c0007", -- 15668
		x"15400015", -- 1566c
		x"46001540", -- 15670
		x"00154600", -- 15674
		x"51cbfff2", -- 15678
		x"363c000f", -- 1567c
		x"142a0015", -- 15680
		x"b4006618", -- 15684
		x"53034600", -- 15688
		x"142a0015", -- 1568c
		x"b400660c", -- 15690
		x"460051cb", -- 15694
		x"ffe84cdf", -- 15698
		x"000f4e75", -- 1569c
		x"50ed0001", -- 156a0
		x"60f408ea", -- 156a4
		x"00020003", -- 156a8
		x"50ed0000", -- 156ac
		x"4e7508aa", -- 156b0
		x"00020003", -- 156b4
		x"422d0000", -- 156b8
		x"4e7548e7", -- 156bc
		x"c0004280", -- 156c0
		x"34801540", -- 156c4
		x"0017122a", -- 156c8
		x"00030201", -- 156cc
		x"00cf6630", -- 156d0
		x"52004a2a", -- 156d4
		x"00116628", -- 156d8
		x"52004a2a", -- 156dc
		x"00136620", -- 156e0
		x"52004a2a", -- 156e4
		x"00196618", -- 156e8
		x"52004a2a", -- 156ec
		x"001b6610", -- 156f0
		x"52004a2a", -- 156f4
		x"001d6608", -- 156f8
		x"52004a2a", -- 156fc
		x"001f6704", -- 15700
		x"50ed0001", -- 15704
		x"4cdf0003", -- 15708
		x"4e75002a", -- 1570c
		x"00110019", -- 15710
		x"2f3c0000", -- 15714
		x"00784eb9", -- 15718
		x"0000526e", -- 1571c
		x"022a00ee", -- 15720
		x"00194e75", -- 15724
		x"61e4002a", -- 15728
		x"00800019", -- 1572c
		x"157c0040", -- 15730
		x"0017157c", -- 15734
		x"005e0015", -- 15738
		x"157c003e", -- 1573c
		x"0015157c", -- 15740
		x"00000017", -- 15744
		x"4e75284a", -- 15748
		x"4eb90001", -- 1574c
		x"504256ed", -- 15750
		x"00016100", -- 15754
		x"ff664a2d", -- 15758
		x"00016704", -- 1575c
		x"50ed0001", -- 15760
		x"4e750001", -- 15764
		x"4e56fffc", -- 15768
		x"206e0008", -- 1576c
		x"22680008", -- 15770
		x"2d690004", -- 15774
		x"fffc2f2d", -- 15778
		x"fff62f0e", -- 1577c
		x"487a0022", -- 15780
		x"2b4ffff6", -- 15784
		x"226efffc", -- 15788
		x"70001029", -- 1578c
		x"00052140", -- 15790
		x"fffc2b6f", -- 15794
		x"0008fff6", -- 15798
		x"defc000c", -- 1579c
		x"4efa0010", -- 157a0
		x"2c5f2b5f", -- 157a4
		x"fff63b7c", -- 157a8
		x"0045fffe", -- 157ac
		x"4e4a598f", -- 157b0
		x"206e0008", -- 157b4
		x"2f28fffc", -- 157b8
		x"2f2e000c", -- 157bc
		x"4eb90000", -- 157c0
		x"a9d4201f", -- 157c4
		x"b0ae0010", -- 157c8
		x"6700000a", -- 157cc
		x"3b7c0046", -- 157d0
		x"fffe4e4a", -- 157d4
		x"4e5e205f", -- 157d8
		x"defc000c", -- 157dc
		x"4ed00001", -- 157e0
		x"4e56fff0", -- 157e4
		x"206e0008", -- 157e8
		x"22680008", -- 157ec
		x"2d690004", -- 157f0
		x"fff02d7c", -- 157f4
		x"00000004", -- 157f8
		x"fff853ae", -- 157fc
		x"fff82d7c", -- 15800
		x"00000010", -- 15804
		x"fffc53ae", -- 15808
		x"fffc202e", -- 1580c
		x"fff8ed80", -- 15810
		x"d0aefffc", -- 15814
		x"2d40fff4", -- 15818
		x"2f2dfff6", -- 1581c
		x"2f0e487a", -- 15820
		x"001e2b4f", -- 15824
		x"fff6206e", -- 15828
		x"fff0116e", -- 1582c
		x"fff70005", -- 15830
		x"2b6f0008", -- 15834
		x"fff6defc", -- 15838
		x"000c4efa", -- 1583c
		x"00102c5f", -- 15840
		x"2b5ffff6", -- 15844
		x"3b7c0007", -- 15848
		x"fffe4e4a", -- 1584c
		x"2f2efff4", -- 15850
		x"2f3c0000", -- 15854
		x"00cf2f2e", -- 15858
		x"00084eba", -- 1585c
		x"ff080cae", -- 15860
		x"00000000", -- 15864
		x"fffc6e9e", -- 15868
		x"0cae0000", -- 1586c
		x"0000fff8", -- 15870
		x"6e884e5e", -- 15874
		x"2e9f4e75", -- 15878
		x"00014e56", -- 1587c
		x"fffc206e", -- 15880
		x"00082268", -- 15884
		x"00082d69", -- 15888
		x"0004fffc", -- 1588c
		x"2f2dfff6", -- 15890
		x"2f0e487a", -- 15894
		x"001e2b4f", -- 15898
		x"fff6226e", -- 1589c
		x"fffc137c", -- 158a0
		x"ff000023", -- 158a4
		x"2b6f0008", -- 158a8
		x"fff6defc", -- 158ac
		x"000c4efa", -- 158b0
		x"00102c5f", -- 158b4
		x"2b5ffff6", -- 158b8
		x"3b7c000e", -- 158bc
		x"fffe4e4a", -- 158c0
		x"2f2dfff6", -- 158c4
		x"2f0e487a", -- 158c8
		x"001e2b4f", -- 158cc
		x"fff6206e", -- 158d0
		x"fffc117c", -- 158d4
		x"ff010037", -- 158d8
		x"2b6f0008", -- 158dc
		x"fff6defc", -- 158e0
		x"000c4efa", -- 158e4
		x"00102c5f", -- 158e8
		x"2b5ffff6", -- 158ec
		x"3b7c001a", -- 158f0
		x"fffe4e4a", -- 158f4
		x"2f2dfff6", -- 158f8
		x"2f0e487a", -- 158fc
		x"001e2b4f", -- 15900
		x"fff6206e", -- 15904
		x"fffc117c", -- 15908
		x"ff04003d", -- 1590c
		x"2b6f0008", -- 15910
		x"fff6defc", -- 15914
		x"000c4efa", -- 15918
		x"00102c5f", -- 1591c
		x"2b5ffff6", -- 15920
		x"3b7c0023", -- 15924
		x"fffe4e4a", -- 15928
		x"42a72f3c", -- 1592c
		x"000000ff", -- 15930
		x"2f2e0008", -- 15934
		x"4ebafe2e", -- 15938
		x"4e5e2e9f", -- 1593c
		x"4e750001", -- 15940
		x"4e56fff8", -- 15944
		x"2f2e0008", -- 15948
		x"4ebaff30", -- 1594c
		x"206e0008", -- 15950
		x"2d680008", -- 15954
		x"fffc226e", -- 15958
		x"fffc2d69", -- 1595c
		x"0004fff8", -- 15960
		x"2f2dfff6", -- 15964
		x"2f0e487a", -- 15968
		x"001e2b4f", -- 1596c
		x"fff6246e", -- 15970
		x"fff8157c", -- 15974
		x"ff200025", -- 15978
		x"2b6f0008", -- 1597c
		x"fff6defc", -- 15980
		x"000c4efa", -- 15984
		x"00102c5f", -- 15988
		x"2b5ffff6", -- 1598c
		x"3b7c0011", -- 15990
		x"fffe4e4a", -- 15994
		x"2f3c0000", -- 15998
		x"00112f3c", -- 1599c
		x"000000ff", -- 159a0
		x"2f2e0008", -- 159a4
		x"4ebafdbe", -- 159a8
		x"206efffc", -- 159ac
		x"2f280004", -- 159b0
		x"42274eb9", -- 159b4
		x"00016788", -- 159b8
		x"4e5e2e9f", -- 159bc
		x"4e750001", -- 159c0
		x"4e56fff8", -- 159c4
		x"2f2e0008", -- 159c8
		x"4ebafeb0", -- 159cc
		x"206e0008", -- 159d0
		x"2d680008", -- 159d4
		x"fffc226e", -- 159d8
		x"fffc2d69", -- 159dc
		x"0004fff8", -- 159e0
		x"2f2dfff6", -- 159e4
		x"2f0e487a", -- 159e8
		x"00242b4f", -- 159ec
		x"fff6246e", -- 159f0
		x"fff8157c", -- 159f4
		x"ff600025", -- 159f8
		x"157cff20", -- 159fc
		x"00252b6f", -- 15a00
		x"0008fff6", -- 15a04
		x"defc000c", -- 15a08
		x"4efa0010", -- 15a0c
		x"2c5f2b5f", -- 15a10
		x"fff63b7c", -- 15a14
		x"0011fffe", -- 15a18
		x"4e4a2f3c", -- 15a1c
		x"00000031", -- 15a20
		x"2f3c0000", -- 15a24
		x"00ff2f2e", -- 15a28
		x"00084eba", -- 15a2c
		x"fd38206e", -- 15a30
		x"fffc2f28", -- 15a34
		x"00044227", -- 15a38
		x"4eb90001", -- 15a3c
		x"67884e5e", -- 15a40
		x"2e9f4e75", -- 15a44
		x"00014e56", -- 15a48
		x"fffc4a2e", -- 15a4c
		x"000c6700", -- 15a50
		x"000e2d7c", -- 15a54
		x"00000001", -- 15a58
		x"fffc6000", -- 15a5c
		x"000642ae", -- 15a60
		x"fffc2f2d", -- 15a64
		x"fff62f0e", -- 15a68
		x"487a002a", -- 15a6c
		x"2b4ffff6", -- 15a70
		x"206e0008", -- 15a74
		x"22680008", -- 15a78
		x"22690004", -- 15a7c
		x"70001029", -- 15a80
		x"00292140", -- 15a84
		x"fffc2b6f", -- 15a88
		x"0008fff6", -- 15a8c
		x"defc000c", -- 15a90
		x"4efa0010", -- 15a94
		x"2c5f2b5f", -- 15a98
		x"fff63b7c", -- 15a9c
		x"002bfffe", -- 15aa0
		x"4e4a206e", -- 15aa4
		x"00082028", -- 15aa8
		x"fffcb0ae", -- 15aac
		x"fffc6700", -- 15ab0
		x"000a3b7c", -- 15ab4
		x"002cfffe", -- 15ab8
		x"4e4a4e5e", -- 15abc
		x"205f5c4f", -- 15ac0
		x"4ed00001", -- 15ac4
		x"4e56fff8", -- 15ac8
		x"2f2e0008", -- 15acc
		x"4ebafdac", -- 15ad0
		x"206e0008", -- 15ad4
		x"2d680008", -- 15ad8
		x"fffc226e", -- 15adc
		x"fffc2d69", -- 15ae0
		x"0004fff8", -- 15ae4
		x"2f2dfff6", -- 15ae8
		x"2f0e487a", -- 15aec
		x"001e2b4f", -- 15af0
		x"fff6246e", -- 15af4
		x"fff8157c", -- 15af8
		x"ff000037", -- 15afc
		x"2b6f0008", -- 15b00
		x"fff6defc", -- 15b04
		x"000c4efa", -- 15b08
		x"00102c5f", -- 15b0c
		x"2b5ffff6", -- 15b10
		x"3b7c001a", -- 15b14
		x"fffe4e4a", -- 15b18
		x"42272f2e", -- 15b1c
		x"00084eba", -- 15b20
		x"ff262f2d", -- 15b24
		x"fff62f0e", -- 15b28
		x"487a001e", -- 15b2c
		x"2b4ffff6", -- 15b30
		x"206efff8", -- 15b34
		x"117cff20", -- 15b38
		x"00252b6f", -- 15b3c
		x"0008fff6", -- 15b40
		x"defc000c", -- 15b44
		x"4efa0010", -- 15b48
		x"2c5f2b5f", -- 15b4c
		x"fff63b7c", -- 15b50
		x"0011fffe", -- 15b54
		x"4e4a1f3c", -- 15b58
		x"00012f2e", -- 15b5c
		x"00084eba", -- 15b60
		x"fee6206e", -- 15b64
		x"fffc2f28", -- 15b68
		x"00044227", -- 15b6c
		x"4eb90001", -- 15b70
		x"67884e5e", -- 15b74
		x"2e9f4e75", -- 15b78
		x"00004e56", -- 15b7c
		x"fffc206e", -- 15b80
		x"00082f28", -- 15b84
		x"00044227", -- 15b88
		x"4eb90001", -- 15b8c
		x"67882f0e", -- 15b90
		x"4ebafc4e", -- 15b94
		x"2f0e4eba", -- 15b98
		x"fda82f0e", -- 15b9c
		x"4ebafe22", -- 15ba0
		x"2f0e4eba", -- 15ba4
		x"ff204e5e", -- 15ba8
		x"2e9f4e75", -- 15bac
		x"20202020", -- 15bb0
		x"696e7465", -- 15bb4
		x"72666163", -- 15bb8
		x"6520636f", -- 15bbc
		x"6e666967", -- 15bc0
		x"75726174", -- 15bc4
		x"696f6e20", -- 15bc8
		x"6572726f", -- 15bcc
		x"72202020", -- 15bd0
		x"20202020", -- 15bd4
		x"20202020", -- 15bd8
		x"66757365", -- 15bdc
		x"20627572", -- 15be0
		x"6e656420", -- 15be4
		x"6f757420", -- 15be8
		x"20202020", -- 15bec
		x"20202020", -- 15bf0
		x"20202020", -- 15bf4
		x"20202020", -- 15bf8
		x"20202020", -- 15bfc
		x"20202020", -- 15c00
		x"72656769", -- 15c04
		x"73746572", -- 15c08
		x"20746573", -- 15c0c
		x"74206661", -- 15c10
		x"696c6564", -- 15c14
		x"20202020", -- 15c18
		x"20202020", -- 15c1c
		x"20202020", -- 15c20
		x"20202020", -- 15c24
		x"5475726e", -- 15c28
		x"204f4646", -- 15c2c
		x"20414c4c", -- 15c30
		x"20534353", -- 15c34
		x"49206465", -- 15c38
		x"76696365", -- 15c3c
		x"732e2020", -- 15c40
		x"20202020", -- 15c44
		x"20202020", -- 15c48
		x"20202020", -- 15c4c
		x"44697363", -- 15c50
		x"6f6e6e65", -- 15c54
		x"63742063", -- 15c58
		x"61626c65", -- 15c5c
		x"20617420", -- 15c60
		x"6e656172", -- 15c64
		x"65737420", -- 15c68
		x"64657669", -- 15c6c
		x"63652e20", -- 15c70
		x"20202020", -- 15c74
		x"20202020", -- 15c78
		x"6c6f6f70", -- 15c7c
		x"20626163", -- 15c80
		x"6b207465", -- 15c84
		x"73742066", -- 15c88
		x"61696c65", -- 15c8c
		x"64202020", -- 15c90
		x"20202020", -- 15c94
		x"20202020", -- 15c98
		x"20202020", -- 15c9c
		x"41747461", -- 15ca0
		x"63682044", -- 15ca4
		x"49464645", -- 15ca8
		x"52454e54", -- 15cac
		x"49414c20", -- 15cb0
		x"74657374", -- 15cb4
		x"20636f6e", -- 15cb8
		x"6e656374", -- 15cbc
		x"6f722e20", -- 15cc0
		x"20202020", -- 15cc4
		x"41747461", -- 15cc8
		x"63682053", -- 15ccc
		x"494e474c", -- 15cd0
		x"452d454e", -- 15cd4
		x"44454420", -- 15cd8
		x"74657374", -- 15cdc
		x"20636f6e", -- 15ce0
		x"6e656374", -- 15ce4
		x"6f722e20", -- 15ce8
		x"20202020", -- 15cec
		x"52656d6f", -- 15cf0
		x"76652074", -- 15cf4
		x"65737420", -- 15cf8
		x"636f6e6e", -- 15cfc
		x"6563746f", -- 15d00
		x"722e2020", -- 15d04
		x"20202020", -- 15d08
		x"20202020", -- 15d0c
		x"20202020", -- 15d10
		x"20202020", -- 15d14
		x"58206361", -- 15d18
		x"6e63656c", -- 15d1c
		x"732c2052", -- 15d20
		x"45545552", -- 15d24
		x"4e20636f", -- 15d28
		x"6e74696e", -- 15d2c
		x"75657320", -- 15d30
		x"74657374", -- 15d34
		x"696e6720", -- 15d38
		x"20202020", -- 15d3c
		x"20202020", -- 15d40
		x"6361626c", -- 15d44
		x"65207465", -- 15d48
		x"73742066", -- 15d4c
		x"61696c65", -- 15d50
		x"64202020", -- 15d54
		x"20202020", -- 15d58
		x"20202020", -- 15d5c
		x"20202020", -- 15d60
		x"20202020", -- 15d64
		x"436f6e6e", -- 15d68
		x"65637420", -- 15d6c
		x"6361626c", -- 15d70
		x"6520746f", -- 15d74
		x"20646576", -- 15d78
		x"6963652e", -- 15d7c
		x"20202020", -- 15d80
		x"20202020", -- 15d84
		x"20202020", -- 15d88
		x"20202020", -- 15d8c
		x"52657374", -- 15d90
		x"6f726520", -- 15d94
		x"706f7765", -- 15d98
		x"7220746f", -- 15d9c
		x"20646576", -- 15da0
		x"69636573", -- 15da4
		x"2e202020", -- 15da8
		x"20202020", -- 15dac
		x"20202020", -- 15db0
		x"20202020", -- 15db4
		x"52455455", -- 15db8
		x"524e2063", -- 15dbc
		x"6f6e7469", -- 15dc0
		x"6e756573", -- 15dc4
		x"206f7065", -- 15dc8
		x"72617469", -- 15dcc
		x"6f6e7320", -- 15dd0
		x"20202020", -- 15dd4
		x"20202020", -- 15dd8
		x"20202020", -- 15ddc
		x"454e5445", -- 15de0
		x"5220636f", -- 15de4
		x"6e74696e", -- 15de8
		x"75657320", -- 15dec
		x"6f706572", -- 15df0
		x"6174696f", -- 15df4
		x"6e732020", -- 15df8
		x"20202020", -- 15dfc
		x"20202020", -- 15e00
		x"20202020", -- 15e04
		x"58206361", -- 15e08
		x"6e63656c", -- 15e0c
		x"732c2045", -- 15e10
		x"4e544552", -- 15e14
		x"20636f6e", -- 15e18
		x"74696e75", -- 15e1c
		x"65732074", -- 15e20
		x"65737469", -- 15e24
		x"6e672020", -- 15e28
		x"20202020", -- 15e2c
		x"20202020", -- 15e30
		x"74657374", -- 15e34
		x"20686f6f", -- 15e38
		x"6420636f", -- 15e3c
		x"6e6e6563", -- 15e40
		x"74656420", -- 15e44
		x"20202020", -- 15e48
		x"20202020", -- 15e4c
		x"20202020", -- 15e50
		x"20202020", -- 15e54
		x"3a207265", -- 15e58
		x"67697374", -- 15e5c
		x"65722074", -- 15e60
		x"65737473", -- 15e64
		x"20003a20", -- 15e68
		x"6c6f6f70", -- 15e6c
		x"20626163", -- 15e70
		x"6b207465", -- 15e74
		x"73747300", -- 15e78
		x"3a206361", -- 15e7c
		x"626c6520", -- 15e80
		x"74657374", -- 15e84
		x"73202020", -- 15e88
		x"20002020", -- 15e8c
		x"20202020", -- 15e90
		x"20202020", -- 15e94
		x"20202020", -- 15e98
		x"20202000", -- 15e9c
		x"00004e56", -- 15ea0
		x"fff82d6e", -- 15ea4
		x"0008fffc", -- 15ea8
		x"206efffc", -- 15eac
		x"2d680018", -- 15eb0
		x"fff842a8", -- 15eb4
		x"00202010", -- 15eb8
		x"6d0007c0", -- 15ebc
		x"b0bc0000", -- 15ec0
		x"00036e00", -- 15ec4
		x"07b6e380", -- 15ec8
		x"323b0006", -- 15ecc
		x"4efb1002", -- 15ed0
		x"00080162", -- 15ed4
		x"06c40732", -- 15ed8
		x"217c0000", -- 15edc
		x"0021001c", -- 15ee0
		x"2268000c", -- 15ee4
		x"22bc0000", -- 15ee8
		x"00012268", -- 15eec
		x"000c237c", -- 15ef0
		x"00000001", -- 15ef4
		x"00042268", -- 15ef8
		x"000c237c", -- 15efc
		x"00000002", -- 15f00
		x"00082028", -- 15f04
		x"00085380", -- 15f08
		x"6d000118", -- 15f0c
		x"b0bc0000", -- 15f10
		x"00026e00", -- 15f14
		x"010ee380", -- 15f18
		x"323b0006", -- 15f1c
		x"4efb1002", -- 15f20
		x"000600ee", -- 15f24
		x"00ee2268", -- 15f28
		x"000c237c", -- 15f2c
		x"ffffffff", -- 15f30
		x"000c2268", -- 15f34
		x"000c237c", -- 15f38
		x"00000002", -- 15f3c
		x"00102268", -- 15f40
		x"000c237c", -- 15f44
		x"00000003", -- 15f48
		x"00142268", -- 15f4c
		x"000c237c", -- 15f50
		x"00000004", -- 15f54
		x"00182268", -- 15f58
		x"000c237c", -- 15f5c
		x"00000005", -- 15f60
		x"001c2268", -- 15f64
		x"000c237c", -- 15f68
		x"00000006", -- 15f6c
		x"00202268", -- 15f70
		x"000c237c", -- 15f74
		x"ffffffff", -- 15f78
		x"00242268", -- 15f7c
		x"000c237c", -- 15f80
		x"00000003", -- 15f84
		x"00282268", -- 15f88
		x"000c237c", -- 15f8c
		x"00000007", -- 15f90
		x"002c2268", -- 15f94
		x"000c237c", -- 15f98
		x"00000005", -- 15f9c
		x"00302268", -- 15fa0
		x"000c237c", -- 15fa4
		x"00000008", -- 15fa8
		x"00342268", -- 15fac
		x"000c237c", -- 15fb0
		x"ffffffff", -- 15fb4
		x"00382268", -- 15fb8
		x"000c237c", -- 15fbc
		x"00000004", -- 15fc0
		x"003c2268", -- 15fc4
		x"000c237c", -- 15fc8
		x"00000009", -- 15fcc
		x"00402268", -- 15fd0
		x"000c237c", -- 15fd4
		x"0000000a", -- 15fd8
		x"00442268", -- 15fdc
		x"000c237c", -- 15fe0
		x"0000000b", -- 15fe4
		x"00482268", -- 15fe8
		x"000c237c", -- 15fec
		x"0000000c", -- 15ff0
		x"004c2268", -- 15ff4
		x"000c237c", -- 15ff8
		x"0000000d", -- 15ffc
		x"00502268", -- 16000
		x"000c237c", -- 16004
		x"fffffffe", -- 16008
		x"00546000", -- 1600c
		x"0022206e", -- 16010
		x"fffc2268", -- 16014
		x"000c237c", -- 16018
		x"fffffffe", -- 1601c
		x"000c6000", -- 16020
		x"000e206e", -- 16024
		x"fffc217c", -- 16028
		x"00000005", -- 1602c
		x"00206000", -- 16030
		x"0656206e", -- 16034
		x"fff842a8", -- 16038
		x"0006226e", -- 1603c
		x"fffc7001", -- 16040
		x"b0a90008", -- 16044
		x"57c08028", -- 16048
		x"000a7207", -- 1604c
		x"b2a90008", -- 16050
		x"5dc18200", -- 16054
		x"6700053a", -- 16058
		x"20290008", -- 1605c
		x"53806d00", -- 16060
		x"0524b0bc", -- 16064
		x"0000000c", -- 16068
		x"6e00051a", -- 1606c
		x"e380323b", -- 16070
		x"00064efb", -- 16074
		x"1002001a", -- 16078
		x"00680120", -- 1607c
		x"01300140", -- 16080
		x"017a0300", -- 16084
		x"0338040a", -- 16088
		x"0422043a", -- 1608c
		x"04520498", -- 16090
		x"117c1001", -- 16094
		x"000a4228", -- 16098
		x"000b4228", -- 1609c
		x"000c2469", -- 160a0
		x"0004082a", -- 160a4
		x"00050001", -- 160a8
		x"56c04400", -- 160ac
		x"08400000", -- 160b0
		x"02000001", -- 160b4
		x"1080246e", -- 160b8
		x"0008216a", -- 160bc
		x"00180002", -- 160c0
		x"06a80000", -- 160c4
		x"000d0002", -- 160c8
		x"20280002", -- 160cc
		x"02800000", -- 160d0
		x"00037204", -- 160d4
		x"9280d3a8", -- 160d8
		x"00026000", -- 160dc
		x"04b42f2d", -- 160e0
		x"fff62f0e", -- 160e4
		x"487a003c", -- 160e8
		x"2b4ffff6", -- 160ec
		x"206e0008", -- 160f0
		x"2f280004", -- 160f4
		x"1f3c0001", -- 160f8
		x"4eb90001", -- 160fc
		x"67882f2e", -- 16100
		x"00084eb9", -- 16104
		x"0001781c", -- 16108
		x"2f2e0008", -- 1610c
		x"42274eb9", -- 16110
		x"00017c02", -- 16114
		x"2b6f0008", -- 16118
		x"fff6defc", -- 1611c
		x"000c4efa", -- 16120
		x"00722c5f", -- 16124
		x"2b5ffff6", -- 16128
		x"206efff8", -- 1612c
		x"4228000a", -- 16130
		x"226efffc", -- 16134
		x"237cffff", -- 16138
		x"fffc0020", -- 1613c
		x"7003b06d", -- 16140
		x"fffe6600", -- 16144
		x"000e217c", -- 16148
		x"00000001", -- 1614c
		x"00066000", -- 16150
		x"00427009", -- 16154
		x"b06dfffe", -- 16158
		x"66000012", -- 1615c
		x"206efff8", -- 16160
		x"217c0000", -- 16164
		x"00020006", -- 16168
		x"60000028", -- 1616c
		x"700ab06d", -- 16170
		x"fffe6600", -- 16174
		x"0012206e", -- 16178
		x"fff8217c", -- 1617c
		x"00000011", -- 16180
		x"00066000", -- 16184
		x"000e206e", -- 16188
		x"fff8217c", -- 1618c
		x"00000003", -- 16190
		x"00066000", -- 16194
		x"03fc206e", -- 16198
		x"fff8217c", -- 1619c
		x"00000004", -- 161a0
		x"00066000", -- 161a4
		x"03ec206e", -- 161a8
		x"fff8217c", -- 161ac
		x"00000005", -- 161b0
		x"00066000", -- 161b4
		x"03dc206e", -- 161b8
		x"fffc7001", -- 161bc
		x"b0680014", -- 161c0
		x"66000012", -- 161c4
		x"226efff8", -- 161c8
		x"237c0000", -- 161cc
		x"000a0006", -- 161d0
		x"6000000e", -- 161d4
		x"206efff8", -- 161d8
		x"217c0000", -- 161dc
		x"00100006", -- 161e0
		x"206efffc", -- 161e4
		x"217c0000", -- 161e8
		x"00020020", -- 161ec
		x"600003a2", -- 161f0
		x"206efffc", -- 161f4
		x"2268000c", -- 161f8
		x"700db011", -- 161fc
		x"6600011e", -- 16200
		x"2f2dfff6", -- 16204
		x"2f0e487a", -- 16208
		x"00f22b4f", -- 1620c
		x"fff62f2e", -- 16210
		x"00081f3c", -- 16214
		x"00014eb9", -- 16218
		x"00017c02", -- 1621c
		x"206efffc", -- 16220
		x"2f280004", -- 16224
		x"4eb90001", -- 16228
		x"8420206e", -- 1622c
		x"fffc2f28", -- 16230
		x"00041f3c", -- 16234
		x"00013f3c", -- 16238
		x"00014eb9", -- 1623c
		x"00018582", -- 16240
		x"206efffc", -- 16244
		x"2f280004", -- 16248
		x"1f3c0001", -- 1624c
		x"42674eb9", -- 16250
		x"00018582", -- 16254
		x"206efffc", -- 16258
		x"2f280004", -- 1625c
		x"42273f3c", -- 16260
		x"00014eb9", -- 16264
		x"00018582", -- 16268
		x"206efffc", -- 1626c
		x"2f280004", -- 16270
		x"42274267", -- 16274
		x"4eb90001", -- 16278
		x"85822079", -- 1627c
		x"fffffed4", -- 16280
		x"7001b028", -- 16284
		x"033f6400", -- 16288
		x"005a2f2e", -- 1628c
		x"00084227", -- 16290
		x"3f3c0001", -- 16294
		x"4eb90001", -- 16298
		x"865e2f2e", -- 1629c
		x"00084227", -- 162a0
		x"42674eb9", -- 162a4
		x"0001865e", -- 162a8
		x"2079ffff", -- 162ac
		x"fed47003", -- 162b0
		x"b028033f", -- 162b4
		x"53c0206e", -- 162b8
		x"fff8c010", -- 162bc
		x"67000024", -- 162c0
		x"2f2e0008", -- 162c4
		x"1f3c0001", -- 162c8
		x"3f3c0001", -- 162cc
		x"4eb90001", -- 162d0
		x"865e2f2e", -- 162d4
		x"00081f3c", -- 162d8
		x"00014267", -- 162dc
		x"4eb90001", -- 162e0
		x"865e206e", -- 162e4
		x"fff8117c", -- 162e8
		x"ff01000b", -- 162ec
		x"2b6f0008", -- 162f0
		x"fff6defc", -- 162f4
		x"000c4efa", -- 162f8
		x"00202c5f", -- 162fc
		x"2b5ffff6", -- 16300
		x"206efff8", -- 16304
		x"217c0000", -- 16308
		x"00060006", -- 1630c
		x"226efffc", -- 16310
		x"237cffff", -- 16314
		x"fffe0020", -- 16318
		x"60000058", -- 1631c
		x"206efffc", -- 16320
		x"2268000c", -- 16324
		x"7058b011", -- 16328
		x"66000016", -- 1632c
		x"226efff8", -- 16330
		x"4229000a", -- 16334
		x"217c0000", -- 16338
		x"00060020", -- 1633c
		x"60000034", -- 16340
		x"206efffc", -- 16344
		x"217c0000", -- 16348
		x"00030020", -- 1634c
		x"7001b068", -- 16350
		x"00146600", -- 16354
		x"0012226e", -- 16358
		x"fff8237c", -- 1635c
		x"0000000a", -- 16360
		x"00066000", -- 16364
		x"000e206e", -- 16368
		x"fff8217c", -- 1636c
		x"00000010", -- 16370
		x"00066000", -- 16374
		x"021c206e", -- 16378
		x"fffc2268", -- 1637c
		x"00040829", -- 16380
		x"00060001", -- 16384
		x"56c04400", -- 16388
		x"4a006700", -- 1638c
		x"0012226e", -- 16390
		x"fff8237c", -- 16394
		x"00000007", -- 16398
		x"00066000", -- 1639c
		x"000e206e", -- 163a0
		x"fff8217c", -- 163a4
		x"00000008", -- 163a8
		x"00066000", -- 163ac
		x"01e4206e", -- 163b0
		x"fff84a28", -- 163b4
		x"000a6600", -- 163b8
		x"0012226e", -- 163bc
		x"fffc237c", -- 163c0
		x"00000006", -- 163c4
		x"00206000", -- 163c8
		x"00b4206e", -- 163cc
		x"fffc2268", -- 163d0
		x"000c700d", -- 163d4
		x"b0116600", -- 163d8
		x"00522f2d", -- 163dc
		x"fff62f0e", -- 163e0
		x"487a0026", -- 163e4
		x"2b4ffff6", -- 163e8
		x"226efff8", -- 163ec
		x"137cff01", -- 163f0
		x"000c2f2e", -- 163f4
		x"00084eba", -- 163f8
		x"f7822b6f", -- 163fc
		x"0008fff6", -- 16400
		x"defc000c", -- 16404
		x"4efa0020", -- 16408
		x"2c5f2b5f", -- 1640c
		x"fff6206e", -- 16410
		x"fff8217c", -- 16414
		x"0000000b", -- 16418
		x"0006226e", -- 1641c
		x"fffc237c", -- 16420
		x"fffffffd", -- 16424
		x"00206000", -- 16428
		x"0054206e", -- 1642c
		x"fffc2268", -- 16430
		x"000c7058", -- 16434
		x"b0116600", -- 16438
		x"000e217c", -- 1643c
		x"00000006", -- 16440
		x"00206000", -- 16444
		x"0038206e", -- 16448
		x"fffc7001", -- 1644c
		x"b0680014", -- 16450
		x"66000012", -- 16454
		x"226efff8", -- 16458
		x"237c0000", -- 1645c
		x"000a0006", -- 16460
		x"6000000e", -- 16464
		x"206efff8", -- 16468
		x"217c0000", -- 1646c
		x"00100006", -- 16470
		x"206efffc", -- 16474
		x"217c0000", -- 16478
		x"00030020", -- 1647c
		x"60000112", -- 16480
		x"206efff8", -- 16484
		x"4a28000c", -- 16488
		x"6700000a", -- 1648c
		x"217c0000", -- 16490
		x"00090006", -- 16494
		x"600000fa", -- 16498
		x"206efff8", -- 1649c
		x"4a28000b", -- 164a0
		x"6700000a", -- 164a4
		x"217c0000", -- 164a8
		x"000c0006", -- 164ac
		x"600000e2", -- 164b0
		x"206efff8", -- 164b4
		x"4a28000b", -- 164b8
		x"6700000a", -- 164bc
		x"217c0000", -- 164c0
		x"000d0006", -- 164c4
		x"600000ca", -- 164c8
		x"206efff8", -- 164cc
		x"1028000b", -- 164d0
		x"8028000c", -- 164d4
		x"67000034", -- 164d8
		x"226efffc", -- 164dc
		x"7001b069", -- 164e0
		x"00146600", -- 164e4
		x"000e217c", -- 164e8
		x"0000000e", -- 164ec
		x"00066000", -- 164f0
		x"000e206e", -- 164f4
		x"fff8217c", -- 164f8
		x"0000000f", -- 164fc
		x"0006206e", -- 16500
		x"fffc217c", -- 16504
		x"00000002", -- 16508
		x"00206000", -- 1650c
		x"0084206e", -- 16510
		x"fff81028", -- 16514
		x"000b8028", -- 16518
		x"000c6600", -- 1651c
		x"0012226e", -- 16520
		x"fffc237c", -- 16524
		x"00000006", -- 16528
		x"00206000", -- 1652c
		x"0054206e", -- 16530
		x"fffc2268", -- 16534
		x"000c700d", -- 16538
		x"b0116600", -- 1653c
		x"000e217c", -- 16540
		x"00000006", -- 16544
		x"00206000", -- 16548
		x"0038206e", -- 1654c
		x"fffc7001", -- 16550
		x"b0680014", -- 16554
		x"66000012", -- 16558
		x"226efff8", -- 1655c
		x"237c0000", -- 16560
		x"000e0006", -- 16564
		x"6000000e", -- 16568
		x"206efff8", -- 1656c
		x"217c0000", -- 16570
		x"000f0006", -- 16574
		x"206efffc", -- 16578
		x"217c0000", -- 1657c
		x"00030020", -- 16580
		x"6000000e", -- 16584
		x"206efffc", -- 16588
		x"217c0000", -- 1658c
		x"00010020", -- 16590
		x"600000f4", -- 16594
		x"206efffc", -- 16598
		x"42a8001c", -- 1659c
		x"4aa80010", -- 165a0
		x"5ec07204", -- 165a4
		x"b2a80010", -- 165a8
		x"5cc1c200", -- 165ac
		x"67000044", -- 165b0
		x"217c0000", -- 165b4
		x"0011001c", -- 165b8
		x"20280010", -- 165bc
		x"2f002f3c", -- 165c0
		x"00000012", -- 165c4
		x"4eb90000", -- 165c8
		x"81b0201f", -- 165cc
		x"206efffc", -- 165d0
		x"43faf882", -- 165d4
		x"d2fcffee", -- 165d8
		x"2468000c", -- 165dc
		x"43f10800", -- 165e0
		x"4c91191f", -- 165e4
		x"4892191f", -- 165e8
		x"15690010", -- 165ec
		x"00106000", -- 165f0
		x"000e206e", -- 165f4
		x"fffc217c", -- 165f8
		x"00000001", -- 165fc
		x"00206000", -- 16600
		x"0086206e", -- 16604
		x"fffc42a8", -- 16608
		x"001c226e", -- 1660c
		x"fff84aa9", -- 16610
		x"00065ec0", -- 16614
		x"7211b2a9", -- 16618
		x"00065cc1", -- 1661c
		x"c2006700", -- 16620
		x"003e217c", -- 16624
		x"00000028", -- 16628
		x"001c2029", -- 1662c
		x"00062f00", -- 16630
		x"2f3c0000", -- 16634
		x"00284eb9", -- 16638
		x"000081b0", -- 1663c
		x"201f206e", -- 16640
		x"fffc43fa", -- 16644
		x"f568d2fc", -- 16648
		x"ffd82468", -- 1664c
		x"000c43f1", -- 16650
		x"08004cd1", -- 16654
		x"197f48d2", -- 16658
		x"197f6000", -- 1665c
		x"001a206e", -- 16660
		x"fff84aa8", -- 16664
		x"00066700", -- 16668
		x"000e226e", -- 1666c
		x"fffc237c", -- 16670
		x"00000001", -- 16674
		x"00206000", -- 16678
		x"000e206e", -- 1667c
		x"fffc217c", -- 16680
		x"00000005", -- 16684
		x"00204e5e", -- 16688
		x"2e9f4e75", -- 1668c
		x"4e754e75", -- 16690
		x"3b7cfff4", -- 16694
		x"fffe2e6d", -- 16698
		x"fff64e75", -- 1669c
		x"3b7cfffc", -- 166a0
		x"fffe60f2", -- 166a4
		x"3b7cfffb", -- 166a8
		x"fffe60ea", -- 166ac
		x"225f2e1f", -- 166b0
		x"2f094e55", -- 166b4
		x"ffde41ed", -- 166b8
		x"ffde30f8", -- 166bc
		x"ff5820f8", -- 166c0
		x"ff5a30f8", -- 166c4
		x"fffa20f8", -- 166c8
		x"fffc49f8", -- 166cc
		x"ff7620dc", -- 166d0
		x"20dc20dc", -- 166d4
		x"31fc4ef9", -- 166d8
		x"ff5821fc", -- 166dc
		x"0001669a", -- 166e0
		x"ff5a31fc", -- 166e4
		x"4ef9fffa", -- 166e8
		x"21fc0001", -- 166ec
		x"6694fffc", -- 166f0
		x"31fc4ef9", -- 166f4
		x"ff7c21fc", -- 166f8
		x"000166a0", -- 166fc
		x"ff7e31fc", -- 16700
		x"4ef9ff76", -- 16704
		x"21fc0001", -- 16708
		x"66a8ff78", -- 1670c
		x"487a000e", -- 16710
		x"2b4ffff6", -- 16714
		x"2f074eb9", -- 16718
		x"00015ea2", -- 1671c
		x"41edffde", -- 16720
		x"31d8ff58", -- 16724
		x"21d8ff5a", -- 16728
		x"31d8fffa", -- 1672c
		x"21d8fffc", -- 16730
		x"49f8ff76", -- 16734
		x"28d828d8", -- 16738
		x"28d84e5d", -- 1673c
		x"4e7508b8", -- 16740
		x"0005fdcc", -- 16744
		x"2f2c0384", -- 16748
		x"296c0384", -- 1674c
		x"0358297c", -- 16750
		x"000166b0", -- 16754
		x"0384487a", -- 16758
		x"001648e7", -- 1675c
		x"fffe240f", -- 16760
		x"4dfa0018", -- 16764
		x"47ec0340", -- 16768
		x"4ef90000", -- 1676c
		x"7d7a295f", -- 16770
		x"03840838", -- 16774
		x"0005fdcc", -- 16778
		x"4e752e42", -- 1677c
		x"4cdf7fff", -- 16780
		x"60ec0000", -- 16784
		x"4e56fffc", -- 16788
		x"2d6e000a", -- 1678c
		x"fffc2f2d", -- 16790
		x"fff62f0e", -- 16794
		x"487a00d6", -- 16798
		x"2b4ffff6", -- 1679c
		x"206efffc", -- 167a0
		x"117cff00", -- 167a4
		x"00012f2d", -- 167a8
		x"fff62f0e", -- 167ac
		x"487a004a", -- 167b0
		x"2b4ffff6", -- 167b4
		x"117cff00", -- 167b8
		x"00234a2e", -- 167bc
		x"00086700", -- 167c0
		x"0014117c", -- 167c4
		x"00100025", -- 167c8
		x"2f3c0000", -- 167cc
		x"001e4eb9", -- 167d0
		x"0000aa8e", -- 167d4
		x"206efffc", -- 167d8
		x"10280007", -- 167dc
		x"02800000", -- 167e0
		x"00077207", -- 167e4
		x"92801141", -- 167e8
		x"00212b6f", -- 167ec
		x"0008fff6", -- 167f0
		x"defc000c", -- 167f4
		x"4efa0010", -- 167f8
		x"2c5f2b5f", -- 167fc
		x"fff63b7c", -- 16800
		x"000dfffe", -- 16804
		x"4e4a206e", -- 16808
		x"fffc117c", -- 1680c
		x"ffc00023", -- 16810
		x"117cff00", -- 16814
		x"0025117c", -- 16818
		x"ff000027", -- 1681c
		x"117cff00", -- 16820
		x"0031117c", -- 16824
		x"ff000039", -- 16828
		x"117cff00", -- 1682c
		x"003b117c", -- 16830
		x"ff00003d", -- 16834
		x"117cff00", -- 16838
		x"0037117c", -- 1683c
		x"ff00002b", -- 16840
		x"4a2e0008", -- 16844
		x"67000018", -- 16848
		x"4a79ffff", -- 1684c
		x"fdc06700", -- 16850
		x"000e2f3c", -- 16854
		x"004c4b40", -- 16858
		x"4eb90000", -- 1685c
		x"aa8e2b6f", -- 16860
		x"0008fff6", -- 16864
		x"defc000c", -- 16868
		x"4efa001c", -- 1686c
		x"2c5f2b5f", -- 16870
		x"fff6700d", -- 16874
		x"b06dfffe", -- 16878
		x"66000004", -- 1687c
		x"4e4a3b7c", -- 16880
		x"0032fffe", -- 16884
		x"4e4a4e5e", -- 16888
		x"205f5c4f", -- 1688c
		x"4ed00000", -- 16890
		x"4e56fff8", -- 16894
		x"422effff", -- 16898
		x"422efffe", -- 1689c
		x"2d7c0001", -- 168a0
		x"86a0fffa", -- 168a4
		x"486efffa", -- 168a8
		x"4eb90000", -- 168ac
		x"521e2f2d", -- 168b0
		x"fff62f0e", -- 168b4
		x"487a0060", -- 168b8
		x"2b4ffff6", -- 168bc
		x"206e0014", -- 168c0
		x"70001028", -- 168c4
		x"002b3d40", -- 168c8
		x"fff8598f", -- 168cc
		x"302efff8", -- 168d0
		x"48c02f00", -- 168d4
		x"2f2e0010", -- 168d8
		x"4eb90000", -- 168dc
		x"a9d4201f", -- 168e0
		x"b0ae000c", -- 168e4
		x"6600001e", -- 168e8
		x"4a2effff", -- 168ec
		x"6700000c", -- 168f0
		x"1d7c0001", -- 168f4
		x"fffe6000", -- 168f8
		x"00081d7c", -- 168fc
		x"0001ffff", -- 16900
		x"60000006", -- 16904
		x"422effff", -- 16908
		x"2b6f0008", -- 1690c
		x"fff6defc", -- 16910
		x"000c4efa", -- 16914
		x"00102c5f", -- 16918
		x"2b5ffff6", -- 1691c
		x"3b7c0026", -- 16920
		x"fffe4e4a", -- 16924
		x"558f486e", -- 16928
		x"fffa4eb9", -- 1692c
		x"00005258", -- 16930
		x"102effff", -- 16934
		x"08400000", -- 16938
		x"c01f802e", -- 1693c
		x"fffe6700", -- 16940
		x"ff6e4a2e", -- 16944
		x"fffe6600", -- 16948
		x"000a3b6e", -- 1694c
		x"000afffe", -- 16950
		x"4e4a4e5e", -- 16954
		x"205fdefc", -- 16958
		x"00104ed0", -- 1695c
		x"00004e56", -- 16960
		x"fff4422e", -- 16964
		x"ffff2d7c", -- 16968
		x"000186a0", -- 1696c
		x"fffa486e", -- 16970
		x"fffa4eb9", -- 16974
		x"0000521e", -- 16978
		x"2d6e000c", -- 1697c
		x"fff42f2d", -- 16980
		x"fff62f0e", -- 16984
		x"487a0022", -- 16988
		x"2b4ffff6", -- 1698c
		x"206efff4", -- 16990
		x"70001028", -- 16994
		x"00293d40", -- 16998
		x"fff82b6f", -- 1699c
		x"0008fff6", -- 169a0
		x"defc000c", -- 169a4
		x"4efa0010", -- 169a8
		x"2c5f2b5f", -- 169ac
		x"fff63b7c", -- 169b0
		x"002bfffe", -- 169b4
		x"4e4a598f", -- 169b8
		x"302efff8", -- 169bc
		x"48c02f00", -- 169c0
		x"598f2f2e", -- 169c4
		x"00084eb9", -- 169c8
		x"0000a9de", -- 169cc
		x"4eb90000", -- 169d0
		x"a9d44a9f", -- 169d4
		x"66000048", -- 169d8
		x"4a6efff8", -- 169dc
		x"6700003c", -- 169e0
		x"2f2dfff6", -- 169e4
		x"2f0e487a", -- 169e8
		x"00242b4f", -- 169ec
		x"fff6206e", -- 169f0
		x"fff4116e", -- 169f4
		x"fff90029", -- 169f8
		x"1d7cff01", -- 169fc
		x"ffff2b6f", -- 16a00
		x"0008fff6", -- 16a04
		x"defc000c", -- 16a08
		x"4efa0010", -- 16a0c
		x"2c5f2b5f", -- 16a10
		x"fff63b7c", -- 16a14
		x"002afffe", -- 16a18
		x"4e4a6000", -- 16a1c
		x"000a3b7c", -- 16a20
		x"002cfffe", -- 16a24
		x"4e4a558f", -- 16a28
		x"486efffa", -- 16a2c
		x"4eb90000", -- 16a30
		x"5258101f", -- 16a34
		x"802effff", -- 16a38
		x"6700ff3e", -- 16a3c
		x"4a2effff", -- 16a40
		x"6600000a", -- 16a44
		x"3b7c0033", -- 16a48
		x"fffe4e4a", -- 16a4c
		x"4e5e205f", -- 16a50
		x"504f4ed0", -- 16a54
		x"00004e56", -- 16a58
		x"00002f2d", -- 16a5c
		x"fff62f0e", -- 16a60
		x"487a0026", -- 16a64
		x"2b4ffff6", -- 16a68
		x"206e0008", -- 16a6c
		x"10280031", -- 16a70
		x"02800000", -- 16a74
		x"00072d40", -- 16a78
		x"000c2b6f", -- 16a7c
		x"0008fff6", -- 16a80
		x"defc000c", -- 16a84
		x"4efa0010", -- 16a88
		x"2c5f2b5f", -- 16a8c
		x"fff63b7c", -- 16a90
		x"0018fffe", -- 16a94
		x"4e4a4e5e", -- 16a98
		x"2e9f4e75", -- 16a9c
		x"00004e56", -- 16aa0
		x"fffc2f2e", -- 16aa4
		x"000c2f3c", -- 16aa8
		x"00000040", -- 16aac
		x"42a72f3c", -- 16ab0
		x"00000039", -- 16ab4
		x"4ebafdda", -- 16ab8
		x"2f2dfff6", -- 16abc
		x"2f0e487a", -- 16ac0
		x"00342b4f", -- 16ac4
		x"fff62d6e", -- 16ac8
		x"000cfffc", -- 16acc
		x"598f2f2e", -- 16ad0
		x"000c4eba", -- 16ad4
		x"ff825097", -- 16ad8
		x"06970000", -- 16adc
		x"0080206e", -- 16ae0
		x"0008201f", -- 16ae4
		x"30802b6f", -- 16ae8
		x"0008fff6", -- 16aec
		x"defc000c", -- 16af0
		x"4efa0020", -- 16af4
		x"2c5f2b5f", -- 16af8
		x"fff67018", -- 16afc
		x"b06dfffe", -- 16b00
		x"66000008", -- 16b04
		x"4e4a6000", -- 16b08
		x"000a3b7c", -- 16b0c
		x"0032fffe", -- 16b10
		x"4e4a4e5e", -- 16b14
		x"205f504f", -- 16b18
		x"4ed00000", -- 16b1c
		x"4e56fffc", -- 16b20
		x"2f2e000c", -- 16b24
		x"2f3c0000", -- 16b28
		x"00402f3c", -- 16b2c
		x"00000040", -- 16b30
		x"2f3c0000", -- 16b34
		x"00394eba", -- 16b38
		x"fd582f2d", -- 16b3c
		x"fff62f0e", -- 16b40
		x"487a002e", -- 16b44
		x"2b4ffff6", -- 16b48
		x"2d6e000c", -- 16b4c
		x"fffc598f", -- 16b50
		x"2f2e000c", -- 16b54
		x"4ebaff00", -- 16b58
		x"5097206e", -- 16b5c
		x"0008201f", -- 16b60
		x"30802b6f", -- 16b64
		x"0008fff6", -- 16b68
		x"defc000c", -- 16b6c
		x"4efa001c", -- 16b70
		x"2c5f2b5f", -- 16b74
		x"fff67018", -- 16b78
		x"b06dfffe", -- 16b7c
		x"66000004", -- 16b80
		x"4e4a3b7c", -- 16b84
		x"0032fffe", -- 16b88
		x"4e4a4e5e", -- 16b8c
		x"205f504f", -- 16b90
		x"4ed00000", -- 16b94
		x"4e56fffc", -- 16b98
		x"2f2dfff6", -- 16b9c
		x"2f0e487a", -- 16ba0
		x"00222b4f", -- 16ba4
		x"fff6206e", -- 16ba8
		x"000c7000", -- 16bac
		x"1028002d", -- 16bb0
		x"2d40fffc", -- 16bb4
		x"2b6f0008", -- 16bb8
		x"fff6defc", -- 16bbc
		x"000c4efa", -- 16bc0
		x"00102c5f", -- 16bc4
		x"2b5ffff6", -- 16bc8
		x"3b7c0028", -- 16bcc
		x"fffe4e4a", -- 16bd0
		x"598f2f2e", -- 16bd4
		x"fffc2f2e", -- 16bd8
		x"00084eb9", -- 16bdc
		x"0000a9d4", -- 16be0
		x"4a9f56c0", -- 16be4
		x"02000001", -- 16be8
		x"1d400010", -- 16bec
		x"4e5e205f", -- 16bf0
		x"504f4ed0", -- 16bf4
		x"00004e56", -- 16bf8
		x"fff642ae", -- 16bfc
		x"fffc558f", -- 16c00
		x"2f2e0016", -- 16c04
		x"2f3c0000", -- 16c08
		x"00024eba", -- 16c0c
		x"ff881d5f", -- 16c10
		x"fff74a2e", -- 16c14
		x"fff76600", -- 16c18
		x"008a7008", -- 16c1c
		x"b0aefffc", -- 16c20
		x"6c00000a", -- 16c24
		x"3b7c003f", -- 16c28
		x"fffe4e4a", -- 16c2c
		x"4a2e0010", -- 16c30
		x"67000032", -- 16c34
		x"206e000c", -- 16c38
		x"4a106700", -- 16c3c
		x"000c206e", -- 16c40
		x"000c4210", -- 16c44
		x"6000000e", -- 16c48
		x"2f2e0016", -- 16c4c
		x"2f2e0012", -- 16c50
		x"4ebafe4c", -- 16c54
		x"2f2e0016", -- 16c58
		x"2f2e0012", -- 16c5c
		x"4ebafebe", -- 16c60
		x"6000003c", -- 16c64
		x"2f2dfff6", -- 16c68
		x"2f0e487a", -- 16c6c
		x"00242b4f", -- 16c70
		x"fff6202e", -- 16c74
		x"0008d0ae", -- 16c78
		x"fffc206e", -- 16c7c
		x"00161140", -- 16c80
		x"00352b6f", -- 16c84
		x"0008fff6", -- 16c88
		x"defc000c", -- 16c8c
		x"4efa0010", -- 16c90
		x"2c5f2b5f", -- 16c94
		x"fff63b7c", -- 16c98
		x"003bfffe", -- 16c9c
		x"4e4a52ae", -- 16ca0
		x"fffc4a2e", -- 16ca4
		x"fff76700", -- 16ca8
		x"ff564e5e", -- 16cac
		x"205fdefc", -- 16cb0
		x"00124ed0", -- 16cb4
		x"00004e56", -- 16cb8
		x"fff642ae", -- 16cbc
		x"fffc558f", -- 16cc0
		x"2f2e0016", -- 16cc4
		x"2f3c0000", -- 16cc8
		x"00014eba", -- 16ccc
		x"fec81d5f", -- 16cd0
		x"fff74a2e", -- 16cd4
		x"fff76600", -- 16cd8
		x"00887008", -- 16cdc
		x"b0aefffc", -- 16ce0
		x"6c00000a", -- 16ce4
		x"3b7c003e", -- 16ce8
		x"fffe4e4a", -- 16cec
		x"4a2e0010", -- 16cf0
		x"6700003e", -- 16cf4
		x"2f2dfff6", -- 16cf8
		x"2f0e487a", -- 16cfc
		x"00222b4f", -- 16d00
		x"fff6206e", -- 16d04
		x"00167000", -- 16d08
		x"10280035", -- 16d0c
		x"2d40fff8", -- 16d10
		x"2b6f0008", -- 16d14
		x"fff6defc", -- 16d18
		x"000c4efa", -- 16d1c
		x"00102c5f", -- 16d20
		x"2b5ffff6", -- 16d24
		x"3b7c003c", -- 16d28
		x"fffe4e4a", -- 16d2c
		x"6000002e", -- 16d30
		x"206e000c", -- 16d34
		x"4a106700", -- 16d38
		x"000c206e", -- 16d3c
		x"000c4210", -- 16d40
		x"6000000e", -- 16d44
		x"2f2e0016", -- 16d48
		x"2f2e0012", -- 16d4c
		x"4ebafd50", -- 16d50
		x"2f2e0016", -- 16d54
		x"2f2e0012", -- 16d58
		x"4ebafdc2", -- 16d5c
		x"52aefffc", -- 16d60
		x"4a2efff7", -- 16d64
		x"6700ff58", -- 16d68
		x"4e5e205f", -- 16d6c
		x"defc0012", -- 16d70
		x"4ed00000", -- 16d74
		x"4e56fff2", -- 16d78
		x"2d6e0012", -- 16d7c
		x"fff22f2d", -- 16d80
		x"fff62f0e", -- 16d84
		x"487a00ea", -- 16d88
		x"2b4ffff6", -- 16d8c
		x"2f2e000e", -- 16d90
		x"2f3c0001", -- 16d94
		x"00004eb9", -- 16d98
		x"000081a8", -- 16d9c
		x"206efff2", -- 16da0
		x"201f1140", -- 16da4
		x"0039202e", -- 16da8
		x"000e6c06", -- 16dac
		x"d0bc0000", -- 16db0
		x"00ffe080", -- 16db4
		x"02800000", -- 16db8
		x"00ff1140", -- 16dbc
		x"003b202e", -- 16dc0
		x"000e0280", -- 16dc4
		x"000000ff", -- 16dc8
		x"1140003d", -- 16dcc
		x"4a2e0008", -- 16dd0
		x"6700000c", -- 16dd4
		x"117c0080", -- 16dd8
		x"00276000", -- 16ddc
		x"000c206e", -- 16de0
		x"fff2117c", -- 16de4
		x"ff000027", -- 16de8
		x"203c0000", -- 16dec
		x"0080d0ae", -- 16df0
		x"000a206e", -- 16df4
		x"fff21140", -- 16df8
		x"0025422e", -- 16dfc
		x"ffff2d7c", -- 16e00
		x"000186a0", -- 16e04
		x"fffa486e", -- 16e08
		x"fffa4eb9", -- 16e0c
		x"0000521e", -- 16e10
		x"206efff2", -- 16e14
		x"70001028", -- 16e18
		x"002d2d40", -- 16e1c
		x"fff6598f", -- 16e20
		x"2f2efff6", -- 16e24
		x"2f3c0000", -- 16e28
		x"00304eb9", -- 16e2c
		x"0000a9d4", -- 16e30
		x"7030b09f", -- 16e34
		x"66000008", -- 16e38
		x"1d7c0001", -- 16e3c
		x"ffff558f", -- 16e40
		x"486efffa", -- 16e44
		x"4eb90000", -- 16e48
		x"5258101f", -- 16e4c
		x"802effff", -- 16e50
		x"67be4a2e", -- 16e54
		x"ffff6600", -- 16e58
		x"000a3b7c", -- 16e5c
		x"003afffe", -- 16e60
		x"4e4a2b6f", -- 16e64
		x"0008fff6", -- 16e68
		x"defc000c", -- 16e6c
		x"4efa001c", -- 16e70
		x"2c5f2b5f", -- 16e74
		x"fff6703a", -- 16e78
		x"b06dfffe", -- 16e7c
		x"66000004", -- 16e80
		x"4e4a3b7c", -- 16e84
		x"0032fffe", -- 16e88
		x"4e4a4e5e", -- 16e8c
		x"205fdefc", -- 16e90
		x"000e4ed0", -- 16e94
		x"00004e56", -- 16e98
		x"fff62d6e", -- 16e9c
		x"000efff6", -- 16ea0
		x"2f2dfff6", -- 16ea4
		x"2f0e487a", -- 16ea8
		x"00462b4f", -- 16eac
		x"fff6206e", -- 16eb0
		x"fff6117c", -- 16eb4
		x"ff000031", -- 16eb8
		x"117cff00", -- 16ebc
		x"0039117c", -- 16ec0
		x"ff00003b", -- 16ec4
		x"117cff04", -- 16ec8
		x"003d7000", -- 16ecc
		x"10280021", -- 16ed0
		x"3d40fffe", -- 16ed4
		x"116effff", -- 16ed8
		x"0037117c", -- 16edc
		x"ff200025", -- 16ee0
		x"2b6f0008", -- 16ee4
		x"fff6defc", -- 16ee8
		x"000c4efa", -- 16eec
		x"00102c5f", -- 16ef0
		x"2b5ffff6", -- 16ef4
		x"3b7c0032", -- 16ef8
		x"fffe4e4a", -- 16efc
		x"2f2e000e", -- 16f00
		x"2f3c0000", -- 16f04
		x"00192f3c", -- 16f08
		x"00000010", -- 16f0c
		x"2f3c0000", -- 16f10
		x"00344eba", -- 16f14
		x"f97c2f2d", -- 16f18
		x"fff62f0e", -- 16f1c
		x"487a001c", -- 16f20
		x"2b4ffff6", -- 16f24
		x"206e000a", -- 16f28
		x"30bc0008", -- 16f2c
		x"2b6f0008", -- 16f30
		x"fff6defc", -- 16f34
		x"000c4efa", -- 16f38
		x"00102c5f", -- 16f3c
		x"2b5ffff6", -- 16f40
		x"3b7c0032", -- 16f44
		x"fffe4e4a", -- 16f48
		x"2f2e000e", -- 16f4c
		x"2f3c0000", -- 16f50
		x"001042a7", -- 16f54
		x"2f3c0000", -- 16f58
		x"00354eba", -- 16f5c
		x"f9342f2d", -- 16f60
		x"fff62f0e", -- 16f64
		x"487a0020", -- 16f68
		x"2b4ffff6", -- 16f6c
		x"7008d06e", -- 16f70
		x"0008206e", -- 16f74
		x"000a3080", -- 16f78
		x"2b6f0008", -- 16f7c
		x"fff6defc", -- 16f80
		x"000c4efa", -- 16f84
		x"00102c5f", -- 16f88
		x"2b5ffff6", -- 16f8c
		x"3b7c0032", -- 16f90
		x"fffe4e4a", -- 16f94
		x"2f2e000e", -- 16f98
		x"2f3c0000", -- 16f9c
		x"00104eba", -- 16fa0
		x"f9be2d6e", -- 16fa4
		x"000efff6", -- 16fa8
		x"2f2dfff6", -- 16fac
		x"2f0e487a", -- 16fb0
		x"00302b4f", -- 16fb4
		x"fff6206e", -- 16fb8
		x"fff64a28", -- 16fbc
		x"002f6700", -- 16fc0
		x"0008117c", -- 16fc4
		x"00020029", -- 16fc8
		x"206efff6", -- 16fcc
		x"116e0009", -- 16fd0
		x"00312b6f", -- 16fd4
		x"0008fff6", -- 16fd8
		x"defc000c", -- 16fdc
		x"4efa0010", -- 16fe0
		x"2c5f2b5f", -- 16fe4
		x"fff63b7c", -- 16fe8
		x"0032fffe", -- 16fec
		x"4e4a1d7c", -- 16ff0
		x"00010012", -- 16ff4
		x"4e5e205f", -- 16ff8
		x"defc000a", -- 16ffc
		x"4ed00000", -- 17000
		x"4e56ffea", -- 17004
		x"2d7c0000", -- 17008
		x"0008ffee", -- 1700c
		x"598f2f2e", -- 17010
		x"000c4eba", -- 17014
		x"fa422d5f", -- 17018
		x"fff27000", -- 1701c
		x"222effee", -- 17020
		x"53812d41", -- 17024
		x"ffeab0ae", -- 17028
		x"ffea6e00", -- 1702c
		x"01122d40", -- 17030
		x"fff82f2e", -- 17034
		x"000c2f2e", -- 17038
		x"00084eba", -- 1703c
		x"fa62202e", -- 17040
		x"fff2c03c", -- 17044
		x"ff016600", -- 17048
		x"00362f2d", -- 1704c
		x"fff62f0e", -- 17050
		x"487a001e", -- 17054
		x"2b4ffff6", -- 17058
		x"206e000c", -- 1705c
		x"116efffb", -- 17060
		x"00372b6f", -- 17064
		x"0008fff6", -- 17068
		x"defc000c", -- 1706c
		x"4efa0010", -- 17070
		x"2c5f2b5f", -- 17074
		x"fff63b7c", -- 17078
		x"001afffe", -- 1707c
		x"4e4a2f2d", -- 17080
		x"fff62f0e", -- 17084
		x"487a001e", -- 17088
		x"2b4ffff6", -- 1708c
		x"206e000c", -- 17090
		x"117c00e0", -- 17094
		x"00252b6f", -- 17098
		x"0008fff6", -- 1709c
		x"defc000c", -- 170a0
		x"4efa0010", -- 170a4
		x"2c5f2b5f", -- 170a8
		x"fff63b7c", -- 170ac
		x"0011fffe", -- 170b0
		x"4e4a2f2e", -- 170b4
		x"000c2f2e", -- 170b8
		x"00084eba", -- 170bc
		x"fa60082e", -- 170c0
		x"0000fff5", -- 170c4
		x"6700003a", -- 170c8
		x"2f2dfff6", -- 170cc
		x"2f0e487a", -- 170d0
		x"00222b4f", -- 170d4
		x"fff6206e", -- 170d8
		x"000c7000", -- 170dc
		x"10280037", -- 170e0
		x"3d40fff6", -- 170e4
		x"2b6f0008", -- 170e8
		x"fff6defc", -- 170ec
		x"000c4efa", -- 170f0
		x"00102c5f", -- 170f4
		x"2b5ffff6", -- 170f8
		x"3b7c001b", -- 170fc
		x"fffe4e4a", -- 17100
		x"2f2dfff6", -- 17104
		x"2f0e487a", -- 17108
		x"001e2b4f", -- 1710c
		x"fff6206e", -- 17110
		x"000c117c", -- 17114
		x"00c00025", -- 17118
		x"2b6f0008", -- 1711c
		x"fff6defc", -- 17120
		x"000c4efa", -- 17124
		x"00102c5f", -- 17128
		x"2b5ffff6", -- 1712c
		x"3b7c0011", -- 17130
		x"fffe4e4a", -- 17134
		x"202efff8", -- 17138
		x"52806800", -- 1713c
		x"feea4e5e", -- 17140
		x"205f504f", -- 17144
		x"4ed00000", -- 17148
		x"4e56ffec", -- 1714c
		x"598f2f2e", -- 17150
		x"000c4eba", -- 17154
		x"f9022d5f", -- 17158
		x"fff62d7c", -- 1715c
		x"00000008", -- 17160
		x"fff02f2e", -- 17164
		x"000c2f2e", -- 17168
		x"00084eba", -- 1716c
		x"f9321d7c", -- 17170
		x"f901fff5", -- 17174
		x"2f2e000c", -- 17178
		x"2f2efff0", -- 1717c
		x"2f3c0000", -- 17180
		x"00044227", -- 17184
		x"4ebafbee", -- 17188
		x"42aefffc", -- 1718c
		x"202efffc", -- 17190
		x"b0aefff0", -- 17194
		x"6c00004c", -- 17198
		x"2f2e000c", -- 1719c
		x"2f2e0008", -- 171a0
		x"202efff6", -- 171a4
		x"c03cff01", -- 171a8
		x"0200ff01", -- 171ac
		x"1f00486e", -- 171b0
		x"fff52f2e", -- 171b4
		x"fffc4eba", -- 171b8
		x"fa3e2f2e", -- 171bc
		x"000c2f2e", -- 171c0
		x"0008202e", -- 171c4
		x"fff6c03c", -- 171c8
		x"ff010200", -- 171cc
		x"ff011f00", -- 171d0
		x"486efff5", -- 171d4
		x"2f2efffc", -- 171d8
		x"4ebafadc", -- 171dc
		x"50aefffc", -- 171e0
		x"60aa2f2e", -- 171e4
		x"000c2f3c", -- 171e8
		x"00000010", -- 171ec
		x"4ebaf770", -- 171f0
		x"2d6e000c", -- 171f4
		x"ffec2f2d", -- 171f8
		x"fff62f0e", -- 171fc
		x"487a0026", -- 17200
		x"2b4ffff6", -- 17204
		x"206effec", -- 17208
		x"4a28002f", -- 1720c
		x"67000008", -- 17210
		x"117c0002", -- 17214
		x"00292b6f", -- 17218
		x"0008fff6", -- 1721c
		x"defc000c", -- 17220
		x"4efa0010", -- 17224
		x"2c5f2b5f", -- 17228
		x"fff63b7c", -- 1722c
		x"0032fffe", -- 17230
		x"4e4a4e5e", -- 17234
		x"205f504f", -- 17238
		x"4ed00001", -- 1723c
		x"4e56fffc", -- 17240
		x"2f2dfff6", -- 17244
		x"2f0e487a", -- 17248
		x"01762b4f", -- 1724c
		x"fff64aae", -- 17250
		x"000e6600", -- 17254
		x"0012206e", -- 17258
		x"0008217c", -- 1725c
		x"00000010", -- 17260
		x"ffe66000", -- 17264
		x"000e206e", -- 17268
		x"0008217c", -- 1726c
		x"00000020", -- 17270
		x"ffe6206e", -- 17274
		x"00082028", -- 17278
		x"ffe65080", -- 1727c
		x"33c00050", -- 17280
		x"0014202e", -- 17284
		x"000ee180", -- 17288
		x"43f90050", -- 1728c
		x"0000d2fc", -- 17290
		x"010043f1", -- 17294
		x"08002d49", -- 17298
		x"fffc4a28", -- 1729c
		x"000e6700", -- 172a0
		x"00222028", -- 172a4
		x"fff86c02", -- 172a8
		x"5680e480", -- 172ac
		x"5380226e", -- 172b0
		x"fffc2340", -- 172b4
		x"0004217c", -- 172b8
		x"00000100", -- 172bc
		x"ffe66000", -- 172c0
		x"001e206e", -- 172c4
		x"00082028", -- 172c8
		x"fff86c02", -- 172cc
		x"5280e280", -- 172d0
		x"5380226e", -- 172d4
		x"fffc2340", -- 172d8
		x"000442a8", -- 172dc
		x"ffe6206e", -- 172e0
		x"0008226e", -- 172e4
		x"fffc22a8", -- 172e8
		x"00104a2e", -- 172ec
		x"000c6700", -- 172f0
		x"000c2168", -- 172f4
		x"ffe6ffe6", -- 172f8
		x"6000000a", -- 172fc
		x"206e0008", -- 17300
		x"58a8ffe6", -- 17304
		x"206e0008", -- 17308
		x"2028ffe6", -- 1730c
		x"d0bc0000", -- 17310
		x"80005080", -- 17314
		x"5480226e", -- 17318
		x"fffc3340", -- 1731c
		x"00084228", -- 17320
		x"ffee217c", -- 17324
		x"000186a0", -- 17328
		x"ffea4868", -- 1732c
		x"ffea4eb9", -- 17330
		x"0000521e", -- 17334
		x"2f2dfff6", -- 17338
		x"2f0e487a", -- 1733c
		x"00262b4f", -- 17340
		x"fff6206e", -- 17344
		x"fffc226e", -- 17348
		x"00087000", -- 1734c
		x"3028000a", -- 17350
		x"2340ffe6", -- 17354
		x"2b6f0008", -- 17358
		x"fff6defc", -- 1735c
		x"000c4efa", -- 17360
		x"00102c5f", -- 17364
		x"2b5ffff6", -- 17368
		x"3b7c003e", -- 1736c
		x"fffe4e4a", -- 17370
		x"206e0008", -- 17374
		x"08280000", -- 17378
		x"ffe96700", -- 1737c
		x"0008117c", -- 17380
		x"0001ffee", -- 17384
		x"558f206e", -- 17388
		x"00084868", -- 1738c
		x"ffea4eb9", -- 17390
		x"00005258", -- 17394
		x"206e0008", -- 17398
		x"101f8028", -- 1739c
		x"ffee6794", -- 173a0
		x"4a28ffee", -- 173a4
		x"6600000a", -- 173a8
		x"3b7c0041", -- 173ac
		x"fffe4e4a", -- 173b0
		x"2b6f0008", -- 173b4
		x"fff6defc", -- 173b8
		x"000c4efa", -- 173bc
		x"00282c5f", -- 173c0
		x"2b5ffff6", -- 173c4
		x"703eb06d", -- 173c8
		x"fffe57c0", -- 173cc
		x"7241b26d", -- 173d0
		x"fffe57c1", -- 173d4
		x"82006700", -- 173d8
		x"00044e4a", -- 173dc
		x"3b7c0040", -- 173e0
		x"fffe4e4a", -- 173e4
		x"4e5e205f", -- 173e8
		x"defc000a", -- 173ec
		x"4ed00001", -- 173f0
		x"4e560000", -- 173f4
		x"4aae000e", -- 173f8
		x"66000012", -- 173fc
		x"206e0008", -- 17400
		x"217c0000", -- 17404
		x"0001ffe6", -- 17408
		x"6000000e", -- 1740c
		x"206e0008", -- 17410
		x"217c0000", -- 17414
		x"0002ffe6", -- 17418
		x"4a2e000c", -- 1741c
		x"6700000e", -- 17420
		x"206e0008", -- 17424
		x"58a8ffe6", -- 17428
		x"6000000c", -- 1742c
		x"206e0008", -- 17430
		x"2168ffe6", -- 17434
		x"ffe6206e", -- 17438
		x"00084a28", -- 1743c
		x"000e6700", -- 17440
		x"000a50a8", -- 17444
		x"ffe66000", -- 17448
		x"000c206e", -- 1744c
		x"00082168", -- 17450
		x"ffe6ffe6", -- 17454
		x"2f2dfff6", -- 17458
		x"2f0e487a", -- 1745c
		x"00222b4f", -- 17460
		x"fff6206e", -- 17464
		x"0008226e", -- 17468
		x"00121368", -- 1746c
		x"ffe90003", -- 17470
		x"2b6f0008", -- 17474
		x"fff6defc", -- 17478
		x"000c4efa", -- 1747c
		x"00102c5f", -- 17480
		x"2b5ffff6", -- 17484
		x"3b7c0004", -- 17488
		x"fffe4e4a", -- 1748c
		x"4e5e205f", -- 17490
		x"defc000e", -- 17494
		x"4ed00001", -- 17498
		x"4e560000", -- 1749c
		x"2f2dfff6", -- 174a0
		x"2f0e487a", -- 174a4
		x"001e2b4f", -- 174a8
		x"fff6206e", -- 174ac
		x"000c117c", -- 174b0
		x"00000003", -- 174b4
		x"2b6f0008", -- 174b8
		x"fff6defc", -- 174bc
		x"000c4efa", -- 174c0
		x"00102c5f", -- 174c4
		x"2b5ffff6", -- 174c8
		x"3b7c0004", -- 174cc
		x"fffe4e4a", -- 174d0
		x"4e5e205f", -- 174d4
		x"504f4ed0", -- 174d8
		x"00004e56", -- 174dc
		x"ffe22d6e", -- 174e0
		x"0014fffc", -- 174e4
		x"58aefffc", -- 174e8
		x"2d7c0000", -- 174ec
		x"0008fff8", -- 174f0
		x"598f2f2e", -- 174f4
		x"00144eba", -- 174f8
		x"f55e2d5f", -- 174fc
		x"fff47000", -- 17500
		x"222efff8", -- 17504
		x"53812d41", -- 17508
		x"ffe2b0ae", -- 1750c
		x"ffe26e00", -- 17510
		x"001c2d40", -- 17514
		x"fff0206e", -- 17518
		x"0010202e", -- 1751c
		x"fff011ae", -- 17520
		x"fff30800", -- 17524
		x"202efff0", -- 17528
		x"528068de", -- 1752c
		x"2f2e0008", -- 17530
		x"202efff4", -- 17534
		x"c03cff01", -- 17538
		x"0200ff01", -- 1753c
		x"1f002f0e", -- 17540
		x"4ebafcfa", -- 17544
		x"2f2e0014", -- 17548
		x"2f2efffc", -- 1754c
		x"4ebaf550", -- 17550
		x"1d7cf501", -- 17554
		x"ffef2f2e", -- 17558
		x"00142f2e", -- 1755c
		x"fff842a7", -- 17560
		x"1f2e000c", -- 17564
		x"4ebaf80e", -- 17568
		x"082e0000", -- 1756c
		x"fff76700", -- 17570
		x"001e42ae", -- 17574
		x"fff02f2e", -- 17578
		x"00142f2e", -- 1757c
		x"fffc1f3c", -- 17580
		x"ff01486e", -- 17584
		x"ffef2f2e", -- 17588
		x"fff04eba", -- 1758c
		x"f66a2f2e", -- 17590
		x"00142f2e", -- 17594
		x"0008202e", -- 17598
		x"fff4c03c", -- 1759c
		x"ff010200", -- 175a0
		x"ff011f00", -- 175a4
		x"2f0e4eba", -- 175a8
		x"fe48422e", -- 175ac
		x"ffee2d7c", -- 175b0
		x"000186a0", -- 175b4
		x"ffea486e", -- 175b8
		x"ffea4eb9", -- 175bc
		x"0000521e", -- 175c0
		x"2f2dfff6", -- 175c4
		x"2f0e487a", -- 175c8
		x"002e2b4f", -- 175cc
		x"fff6202e", -- 175d0
		x"0008e180", -- 175d4
		x"41f90050", -- 175d8
		x"0000d0fc", -- 175dc
		x"010a7200", -- 175e0
		x"32300800", -- 175e4
		x"2d41ffe6", -- 175e8
		x"2b6f0008", -- 175ec
		x"fff6defc", -- 175f0
		x"000c4efa", -- 175f4
		x"00102c5f", -- 175f8
		x"2b5ffff6", -- 175fc
		x"3b7c0040", -- 17600
		x"fffe4e4a", -- 17604
		x"202effe6", -- 17608
		x"c03cff01", -- 1760c
		x"66000008", -- 17610
		x"1d7c0001", -- 17614
		x"ffee558f", -- 17618
		x"486effea", -- 1761c
		x"4eb90000", -- 17620
		x"5258101f", -- 17624
		x"802effee", -- 17628
		x"67962f2e", -- 1762c
		x"00142f0e", -- 17630
		x"4ebafe66", -- 17634
		x"598f2f2e", -- 17638
		x"ffe62f3c", -- 1763c
		x"0000007f", -- 17640
		x"4eb90000", -- 17644
		x"a9d44a9f", -- 17648
		x"6700000a", -- 1764c
		x"3b7c0042", -- 17650
		x"fffe4e4a", -- 17654
		x"202efff4", -- 17658
		x"c03cff01", -- 1765c
		x"66000018", -- 17660
		x"2f2e0014", -- 17664
		x"2f2efffc", -- 17668
		x"4227486e", -- 1766c
		x"ffef2f2e", -- 17670
		x"fff04eba", -- 17674
		x"f6422f2e", -- 17678
		x"00142f3c", -- 1767c
		x"00000010", -- 17680
		x"4ebaf2dc", -- 17684
		x"2d6e0014", -- 17688
		x"ffe22f2d", -- 1768c
		x"fff62f0e", -- 17690
		x"487a0026", -- 17694
		x"2b4ffff6", -- 17698
		x"206effe2", -- 1769c
		x"4a28002f", -- 176a0
		x"67000008", -- 176a4
		x"117c0002", -- 176a8
		x"00292b6f", -- 176ac
		x"0008fff6", -- 176b0
		x"defc000c", -- 176b4
		x"4efa0010", -- 176b8
		x"2c5f2b5f", -- 176bc
		x"fff63b7c", -- 176c0
		x"0032fffe", -- 176c4
		x"4e4a4e5e", -- 176c8
		x"205fdefc", -- 176cc
		x"00104ed0", -- 176d0
		x"00004e56", -- 176d4
		x"fff62f2d", -- 176d8
		x"fff62f0e", -- 176dc
		x"487a001a", -- 176e0
		x"2b4ffff6", -- 176e4
		x"206e0008", -- 176e8
		x"42502b6f", -- 176ec
		x"0008fff6", -- 176f0
		x"defc000c", -- 176f4
		x"4efa0010", -- 176f8
		x"2c5f2b5f", -- 176fc
		x"fff63b7c", -- 17700
		x"0032fffe", -- 17704
		x"4e4a2f2e", -- 17708
		x"000c2f3c", -- 1770c
		x"00000020", -- 17710
		x"4ebaf24c", -- 17714
		x"2d6e000c", -- 17718
		x"fff62f2d", -- 1771c
		x"fff62f0e", -- 17720
		x"487a0026", -- 17724
		x"2b4ffff6", -- 17728
		x"206efff6", -- 1772c
		x"4a28002f", -- 17730
		x"67000008", -- 17734
		x"117c0002", -- 17738
		x"00292b6f", -- 1773c
		x"0008fff6", -- 17740
		x"defc000c", -- 17744
		x"4efa0010", -- 17748
		x"2c5f2b5f", -- 1774c
		x"fff63b7c", -- 17750
		x"0032fffe", -- 17754
		x"4e4a4e5e", -- 17758
		x"205f504f", -- 1775c
		x"4ed04e75", -- 17760
		x"00014e56", -- 17764
		x"fffc206e", -- 17768
		x"00082268", -- 1776c
		x"00082d69", -- 17770
		x"0004fffc", -- 17774
		x"2f2dfff6", -- 17778
		x"2f0e487a", -- 1777c
		x"001e2b4f", -- 17780
		x"fff6226e", -- 17784
		x"fffc136e", -- 17788
		x"00130003", -- 1778c
		x"2b6f0008", -- 17790
		x"fff6defc", -- 17794
		x"000c4efa", -- 17798
		x"00102c5f", -- 1779c
		x"2b5ffff6", -- 177a0
		x"3b7c0004", -- 177a4
		x"fffe4e4a", -- 177a8
		x"2f2dfff6", -- 177ac
		x"2f0e487a", -- 177b0
		x"00422b4f", -- 177b4
		x"fff6598f", -- 177b8
		x"206efffc", -- 177bc
		x"70001028", -- 177c0
		x"00032f00", -- 177c4
		x"226e0008", -- 177c8
		x"2f29fffc", -- 177cc
		x"4eb90000", -- 177d0
		x"a9d4201f", -- 177d4
		x"b0ae000c", -- 177d8
		x"6700000a", -- 177dc
		x"3b7c0006", -- 177e0
		x"fffe4e4a", -- 177e4
		x"2b6f0008", -- 177e8
		x"fff6defc", -- 177ec
		x"000c4efa", -- 177f0
		x"001c2c5f", -- 177f4
		x"2b5ffff6", -- 177f8
		x"7006b06d", -- 177fc
		x"fffe6600", -- 17800
		x"00044e4a", -- 17804
		x"3b7c0005", -- 17808
		x"fffe4e4a", -- 1780c
		x"4e5e205f", -- 17810
		x"defc000c", -- 17814
		x"4ed00000", -- 17818
		x"4e56fff0", -- 1781c
		x"2d6e0008", -- 17820
		x"fff8206e", -- 17824
		x"fff82d68", -- 17828
		x"0004fff4", -- 1782c
		x"2d680018", -- 17830
		x"fff02f28", -- 17834
		x"00044227", -- 17838
		x"4eb90001", -- 1783c
		x"6788206e", -- 17840
		x"fff04a10", -- 17844
		x"6700000e", -- 17848
		x"2d7c0000", -- 1784c
		x"00cffffc", -- 17850
		x"6000000a", -- 17854
		x"2d7c0000", -- 17858
		x"00c7fffc", -- 1785c
		x"206efff0", -- 17860
		x"4a106700", -- 17864
		x"00182f3c", -- 17868
		x"0000007f", -- 1786c
		x"2f3c0000", -- 17870
		x"000f2f0e", -- 17874
		x"4ebafeec", -- 17878
		x"60000014", -- 1787c
		x"2f3c0000", -- 17880
		x"007f2f3c", -- 17884
		x"00000007", -- 17888
		x"2f0e4eba", -- 1788c
		x"fed642a7", -- 17890
		x"42a72f0e", -- 17894
		x"4ebafecc", -- 17898
		x"206efff0", -- 1789c
		x"4a106700", -- 178a0
		x"00182f3c", -- 178a4
		x"0000007f", -- 178a8
		x"2f3c0000", -- 178ac
		x"000f2f0e", -- 178b0
		x"4ebafeb0", -- 178b4
		x"60000014", -- 178b8
		x"2f3c0000", -- 178bc
		x"007f2f3c", -- 178c0
		x"00000007", -- 178c4
		x"2f0e4eba", -- 178c8
		x"fe9a2f2d", -- 178cc
		x"fff62f0e", -- 178d0
		x"487a001e", -- 178d4
		x"2b4ffff6", -- 178d8
		x"206efff4", -- 178dc
		x"117cff00", -- 178e0
		x"00052b6f", -- 178e4
		x"0008fff6", -- 178e8
		x"defc000c", -- 178ec
		x"4efa0010", -- 178f0
		x"2c5f2b5f", -- 178f4
		x"fff63b7c", -- 178f8
		x"0007fffe", -- 178fc
		x"4e4a2f2d", -- 17900
		x"fff62f0e", -- 17904
		x"487a004c", -- 17908
		x"2b4ffff6", -- 1790c
		x"206efff4", -- 17910
		x"08280007", -- 17914
		x"000756c0", -- 17918
		x"44004a00", -- 1791c
		x"6600000a", -- 17920
		x"3b7c0009", -- 17924
		x"fffe4e4a", -- 17928
		x"206efff4", -- 1792c
		x"08280004", -- 17930
		x"000756c0", -- 17934
		x"44004a00", -- 17938
		x"6700000a", -- 1793c
		x"3b7c0003", -- 17940
		x"fffe4e4a", -- 17944
		x"2b6f0008", -- 17948
		x"fff6defc", -- 1794c
		x"000c4efa", -- 17950
		x"00282c5f", -- 17954
		x"2b5ffff6", -- 17958
		x"7009b06d", -- 1795c
		x"fffe57c0", -- 17960
		x"7203b26d", -- 17964
		x"fffe57c1", -- 17968
		x"82006700", -- 1796c
		x"00044e4a", -- 17970
		x"3b7c0008", -- 17974
		x"fffe4e4a", -- 17978
		x"2f2dfff6", -- 1797c
		x"2f0e487a", -- 17980
		x"001e2b4f", -- 17984
		x"fff6206e", -- 17988
		x"fff4117c", -- 1798c
		x"ff000001", -- 17990
		x"2b6f0008", -- 17994
		x"fff6defc", -- 17998
		x"000c4efa", -- 1799c
		x"00102c5f", -- 179a0
		x"2b5ffff6", -- 179a4
		x"3b7c0001", -- 179a8
		x"fffe4e4a", -- 179ac
		x"2f2dfff6", -- 179b0
		x"2f0e487a", -- 179b4
		x"003c2b4f", -- 179b8
		x"fff6598f", -- 179bc
		x"206efff4", -- 179c0
		x"70001028", -- 179c4
		x"00032f00", -- 179c8
		x"2f3c0000", -- 179cc
		x"00cf4eb9", -- 179d0
		x"0000a9d4", -- 179d4
		x"4a9f6700", -- 179d8
		x"000a3b7c", -- 179dc
		x"0006fffe", -- 179e0
		x"4e4a2b6f", -- 179e4
		x"0008fff6", -- 179e8
		x"defc000c", -- 179ec
		x"4efa001c", -- 179f0
		x"2c5f2b5f", -- 179f4
		x"fff67006", -- 179f8
		x"b06dfffe", -- 179fc
		x"66000004", -- 17a00
		x"4e4a3b7c", -- 17a04
		x"0005fffe", -- 17a08
		x"4e4a206e", -- 17a0c
		x"fff4117c", -- 17a10
		x"ff000005", -- 17a14
		x"4a280005", -- 17a18
		x"66000018", -- 17a1c
		x"117c00ff", -- 17a20
		x"00054a28", -- 17a24
		x"00056700", -- 17a28
		x"000a3b7c", -- 17a2c
		x"000afffe", -- 17a30
		x"4e4a4e5e", -- 17a34
		x"2e9f4e75", -- 17a38
		x"00014e56", -- 17a3c
		x"00002f2d", -- 17a40
		x"fff62f0e", -- 17a44
		x"487a0036", -- 17a48
		x"2b4ffff6", -- 17a4c
		x"206e0008", -- 17a50
		x"2268000a", -- 17a54
		x"22690004", -- 17a58
		x"70001029", -- 17a5c
		x"0023b0ae", -- 17a60
		x"000c6700", -- 17a64
		x"000a3b7c", -- 17a68
		x"0010fffe", -- 17a6c
		x"4e4a2b6f", -- 17a70
		x"0008fff6", -- 17a74
		x"defc000c", -- 17a78
		x"4efa001c", -- 17a7c
		x"2c5f2b5f", -- 17a80
		x"fff67010", -- 17a84
		x"b06dfffe", -- 17a88
		x"66000004", -- 17a8c
		x"4e4a3b7c", -- 17a90
		x"000ffffe", -- 17a94
		x"4e4a4e5e", -- 17a98
		x"205f504f", -- 17a9c
		x"4ed00001", -- 17aa0
		x"4e56fffc", -- 17aa4
		x"206e0008", -- 17aa8
		x"2268000a", -- 17aac
		x"2d690004", -- 17ab0
		x"fffc2f2d", -- 17ab4
		x"fff62f0e", -- 17ab8
		x"487a001e", -- 17abc
		x"2b4ffff6", -- 17ac0
		x"226efffc", -- 17ac4
		x"136e000f", -- 17ac8
		x"00312b6f", -- 17acc
		x"0008fff6", -- 17ad0
		x"defc000c", -- 17ad4
		x"4efa0010", -- 17ad8
		x"2c5f2b5f", -- 17adc
		x"fff63b7c", -- 17ae0
		x"0017fffe", -- 17ae4
		x"4e4a2f2d", -- 17ae8
		x"fff62f0e", -- 17aec
		x"487a002e", -- 17af0
		x"2b4ffff6", -- 17af4
		x"206efffc", -- 17af8
		x"70001028", -- 17afc
		x"0031b0ae", -- 17b00
		x"000c6700", -- 17b04
		x"000a3b7c", -- 17b08
		x"0019fffe", -- 17b0c
		x"4e4a2b6f", -- 17b10
		x"0008fff6", -- 17b14
		x"defc000c", -- 17b18
		x"4efa001c", -- 17b1c
		x"2c5f2b5f", -- 17b20
		x"fff67019", -- 17b24
		x"b06dfffe", -- 17b28
		x"66000004", -- 17b2c
		x"4e4a3b7c", -- 17b30
		x"0018fffe", -- 17b34
		x"4e4a4e5e", -- 17b38
		x"205f504f", -- 17b3c
		x"4ed00001", -- 17b40
		x"4e56fff8", -- 17b44
		x"206e0008", -- 17b48
		x"2d68000a", -- 17b4c
		x"fffc226e", -- 17b50
		x"fffc2d69", -- 17b54
		x"0004fff8", -- 17b58
		x"2f290004", -- 17b5c
		x"42274eb9", -- 17b60
		x"00016788", -- 17b64
		x"2f2dfff6", -- 17b68
		x"2f0e487a", -- 17b6c
		x"00242b4f", -- 17b70
		x"fff6206e", -- 17b74
		x"fff8117c", -- 17b78
		x"ff800031", -- 17b7c
		x"117cff01", -- 17b80
		x"00232b6f", -- 17b84
		x"0008fff6", -- 17b88
		x"defc000c", -- 17b8c
		x"4efa0010", -- 17b90
		x"2c5f2b5f", -- 17b94
		x"fff63b7c", -- 17b98
		x"0017fffe", -- 17b9c
		x"4e4a206e", -- 17ba0
		x"fffc2f28", -- 17ba4
		x"00042f3c", -- 17ba8
		x"00000020", -- 17bac
		x"4eb90001", -- 17bb0
		x"69622f2d", -- 17bb4
		x"fff62f0e", -- 17bb8
		x"487a001e", -- 17bbc
		x"2b4ffff6", -- 17bc0
		x"206efff8", -- 17bc4
		x"117cff00", -- 17bc8
		x"00312b6f", -- 17bcc
		x"0008fff6", -- 17bd0
		x"defc000c", -- 17bd4
		x"4efa0010", -- 17bd8
		x"2c5f2b5f", -- 17bdc
		x"fff63b7c", -- 17be0
		x"0032fffe", -- 17be4
		x"4e4a206e", -- 17be8
		x"fffc2f28", -- 17bec
		x"00044227", -- 17bf0
		x"4eb90001", -- 17bf4
		x"67884e5e", -- 17bf8
		x"2e9f4e75", -- 17bfc
		x"00004e56", -- 17c00
		x"fff02d6e", -- 17c04
		x"000afff4", -- 17c08
		x"206efff4", -- 17c0c
		x"2d680004", -- 17c10
		x"fff02f28", -- 17c14
		x"00044227", -- 17c18
		x"4eb90001", -- 17c1c
		x"67882d7c", -- 17c20
		x"00000001", -- 17c24
		x"fffc2d7c", -- 17c28
		x"ffffffff", -- 17c2c
		x"fff852ae", -- 17c30
		x"fff82f2d", -- 17c34
		x"fff62f0e", -- 17c38
		x"487a001e", -- 17c3c
		x"2b4ffff6", -- 17c40
		x"206efff0", -- 17c44
		x"116efffb", -- 17c48
		x"00212b6f", -- 17c4c
		x"0008fff6", -- 17c50
		x"defc000c", -- 17c54
		x"4efa0010", -- 17c58
		x"2c5f2b5f", -- 17c5c
		x"fff63b7c", -- 17c60
		x"000afffe", -- 17c64
		x"4e4a2f2d", -- 17c68
		x"fff62f0e", -- 17c6c
		x"487a002e", -- 17c70
		x"2b4ffff6", -- 17c74
		x"206efff0", -- 17c78
		x"70001028", -- 17c7c
		x"0021b0ae", -- 17c80
		x"fffc6700", -- 17c84
		x"000a3b7c", -- 17c88
		x"000cfffe", -- 17c8c
		x"4e4a2b6f", -- 17c90
		x"0008fff6", -- 17c94
		x"defc000c", -- 17c98
		x"4efa001c", -- 17c9c
		x"2c5f2b5f", -- 17ca0
		x"fff6700c", -- 17ca4
		x"b06dfffe", -- 17ca8
		x"66000004", -- 17cac
		x"4e4a3b7c", -- 17cb0
		x"000bfffe", -- 17cb4
		x"4e4a202e", -- 17cb8
		x"fffce380", -- 17cbc
		x"2d40fffc", -- 17cc0
		x"0cae0000", -- 17cc4
		x"0007fff8", -- 17cc8
		x"6d00ff64", -- 17ccc
		x"2d7c0000", -- 17cd0
		x"007ffff8", -- 17cd4
		x"52aefff8", -- 17cd8
		x"2f2dfff6", -- 17cdc
		x"2f0e487a", -- 17ce0
		x"001e2b4f", -- 17ce4
		x"fff6206e", -- 17ce8
		x"fff0116e", -- 17cec
		x"fffb0023", -- 17cf0
		x"2b6f0008", -- 17cf4
		x"fff6defc", -- 17cf8
		x"000c4efa", -- 17cfc
		x"00102c5f", -- 17d00
		x"2b5ffff6", -- 17d04
		x"3b7c000e", -- 17d08
		x"fffe4e4a", -- 17d0c
		x"0cae0000", -- 17d10
		x"00fffff8", -- 17d14
		x"6dbe2f2e", -- 17d18
		x"fff82f0e", -- 17d1c
		x"4ebafd1c", -- 17d20
		x"2f2dfff6", -- 17d24
		x"2f0e487a", -- 17d28
		x"001e2b4f", -- 17d2c
		x"fff6206e", -- 17d30
		x"fff0117c", -- 17d34
		x"ff7f0023", -- 17d38
		x"2b6f0008", -- 17d3c
		x"fff6defc", -- 17d40
		x"000c4efa", -- 17d44
		x"00102c5f", -- 17d48
		x"2b5ffff6", -- 17d4c
		x"3b7c000e", -- 17d50
		x"fffe4e4a", -- 17d54
		x"2f3c0000", -- 17d58
		x"007f2f0e", -- 17d5c
		x"4ebafcdc", -- 17d60
		x"2f2dfff6", -- 17d64
		x"2f0e487a", -- 17d68
		x"001e2b4f", -- 17d6c
		x"fff6206e", -- 17d70
		x"fff0117c", -- 17d74
		x"ff000001", -- 17d78
		x"2b6f0008", -- 17d7c
		x"fff6defc", -- 17d80
		x"000c4efa", -- 17d84
		x"00102c5f", -- 17d88
		x"2b5ffff6", -- 17d8c
		x"3b7c0001", -- 17d90
		x"fffe4e4a", -- 17d94
		x"2f3c0000", -- 17d98
		x"00802f0e", -- 17d9c
		x"4ebafc9c", -- 17da0
		x"2d7c0000", -- 17da4
		x"0100fff8", -- 17da8
		x"53aefff8", -- 17dac
		x"598f2f2e", -- 17db0
		x"fff82f3c", -- 17db4
		x"00000012", -- 17db8
		x"4eb90000", -- 17dbc
		x"a9d44a9f", -- 17dc0
		x"66000036", -- 17dc4
		x"2f2dfff6", -- 17dc8
		x"2f0e487a", -- 17dcc
		x"001e2b4f", -- 17dd0
		x"fff6206e", -- 17dd4
		x"fff0116e", -- 17dd8
		x"fffb0025", -- 17ddc
		x"2b6f0008", -- 17de0
		x"fff6defc", -- 17de4
		x"000c4efa", -- 17de8
		x"00102c5f", -- 17dec
		x"2b5ffff6", -- 17df0
		x"3b7c0011", -- 17df4
		x"fffe4e4a", -- 17df8
		x"0cae0000", -- 17dfc
		x"0000fff8", -- 17e00
		x"6ea62f2d", -- 17e04
		x"fff62f0e", -- 17e08
		x"487a002e", -- 17e0c
		x"2b4ffff6", -- 17e10
		x"206efff0", -- 17e14
		x"70001028", -- 17e18
		x"0025b0ae", -- 17e1c
		x"fff86700", -- 17e20
		x"000a3b7c", -- 17e24
		x"0013fffe", -- 17e28
		x"4e4a2b6f", -- 17e2c
		x"0008fff6", -- 17e30
		x"defc000c", -- 17e34
		x"4efa001c", -- 17e38
		x"2c5f2b5f", -- 17e3c
		x"fff67013", -- 17e40
		x"b06dfffe", -- 17e44
		x"66000004", -- 17e48
		x"4e4a3b7c", -- 17e4c
		x"0012fffe", -- 17e50
		x"4e4a2d7c", -- 17e54
		x"00000040", -- 17e58
		x"fff853ae", -- 17e5c
		x"fff82f2d", -- 17e60
		x"fff62f0e", -- 17e64
		x"487a0022", -- 17e68
		x"2b4ffff6", -- 17e6c
		x"202efff8", -- 17e70
		x"e580206e", -- 17e74
		x"fff01140", -- 17e78
		x"00272b6f", -- 17e7c
		x"0008fff6", -- 17e80
		x"defc000c", -- 17e84
		x"4efa0010", -- 17e88
		x"2c5f2b5f", -- 17e8c
		x"fff63b7c", -- 17e90
		x"0014fffe", -- 17e94
		x"4e4a0cae", -- 17e98
		x"00000000", -- 17e9c
		x"fff86eba", -- 17ea0
		x"2f2dfff6", -- 17ea4
		x"2f0e487a", -- 17ea8
		x"00322b4f", -- 17eac
		x"fff6202e", -- 17eb0
		x"fff8e580", -- 17eb4
		x"206efff0", -- 17eb8
		x"72001228", -- 17ebc
		x"0027b081", -- 17ec0
		x"6700000a", -- 17ec4
		x"3b7c0016", -- 17ec8
		x"fffe4e4a", -- 17ecc
		x"2b6f0008", -- 17ed0
		x"fff6defc", -- 17ed4
		x"000c4efa", -- 17ed8
		x"001c2c5f", -- 17edc
		x"2b5ffff6", -- 17ee0
		x"7016b06d", -- 17ee4
		x"fffe6600", -- 17ee8
		x"00044e4a", -- 17eec
		x"3b7c0015", -- 17ef0
		x"fffe4e4a", -- 17ef4
		x"2d7c0000", -- 17ef8
		x"0088fff8", -- 17efc
		x"53aefff8", -- 17f00
		x"2f2efff8", -- 17f04
		x"2f0e4eba", -- 17f08
		x"fb980cae", -- 17f0c
		x"00000080", -- 17f10
		x"fff86ee8", -- 17f14
		x"2d7c0000", -- 17f18
		x"0008fff8", -- 17f1c
		x"53aefff8", -- 17f20
		x"2f2efff8", -- 17f24
		x"2f0e4eba", -- 17f28
		x"fb780cae", -- 17f2c
		x"00000000", -- 17f30
		x"fff86ee8", -- 17f34
		x"2f2dfff6", -- 17f38
		x"2f0e487a", -- 17f3c
		x"001e2b4f", -- 17f40
		x"fff6206e", -- 17f44
		x"fff0117c", -- 17f48
		x"ff000037", -- 17f4c
		x"2b6f0008", -- 17f50
		x"fff6defc", -- 17f54
		x"000c4efa", -- 17f58
		x"00102c5f", -- 17f5c
		x"2b5ffff6", -- 17f60
		x"3b7c001a", -- 17f64
		x"fffe4e4a", -- 17f68
		x"2d7c0000", -- 17f6c
		x"0100fff8", -- 17f70
		x"53aefff8", -- 17f74
		x"2f2dfff6", -- 17f78
		x"2f0e487a", -- 17f7c
		x"001e2b4f", -- 17f80
		x"fff6206e", -- 17f84
		x"fff0116e", -- 17f88
		x"fffb0039", -- 17f8c
		x"2b6f0008", -- 17f90
		x"fff6defc", -- 17f94
		x"000c4efa", -- 17f98
		x"00102c5f", -- 17f9c
		x"2b5ffff6", -- 17fa0
		x"3b7c001d", -- 17fa4
		x"fffe4e4a", -- 17fa8
		x"2f2dfff6", -- 17fac
		x"2f0e487a", -- 17fb0
		x"002e2b4f", -- 17fb4
		x"fff6206e", -- 17fb8
		x"fff07000", -- 17fbc
		x"10280039", -- 17fc0
		x"b0aefff8", -- 17fc4
		x"6700000a", -- 17fc8
		x"3b7c001f", -- 17fcc
		x"fffe4e4a", -- 17fd0
		x"2b6f0008", -- 17fd4
		x"fff6defc", -- 17fd8
		x"000c4efa", -- 17fdc
		x"001c2c5f", -- 17fe0
		x"2b5ffff6", -- 17fe4
		x"701fb06d", -- 17fe8
		x"fffe6600", -- 17fec
		x"00044e4a", -- 17ff0
		x"3b7c001e", -- 17ff4
		x"fffe4e4a", -- 17ff8
		x"0cae0000", -- 17ffc
		x"0000fff8", -- 18000
		x"6e00ff6e", -- 18004
		x"2d7c0000", -- 18008
		x"0100fff8", -- 1800c
		x"53aefff8", -- 18010
		x"2f2dfff6", -- 18014
		x"2f0e487a", -- 18018
		x"001e2b4f", -- 1801c
		x"fff6206e", -- 18020
		x"fff0116e", -- 18024
		x"fffb003b", -- 18028
		x"2b6f0008", -- 1802c
		x"fff6defc", -- 18030
		x"000c4efa", -- 18034
		x"00102c5f", -- 18038
		x"2b5ffff6", -- 1803c
		x"3b7c0020", -- 18040
		x"fffe4e4a", -- 18044
		x"2f2dfff6", -- 18048
		x"2f0e487a", -- 1804c
		x"002e2b4f", -- 18050
		x"fff6206e", -- 18054
		x"fff07000", -- 18058
		x"1028003b", -- 1805c
		x"b0aefff8", -- 18060
		x"6700000a", -- 18064
		x"3b7c0022", -- 18068
		x"fffe4e4a", -- 1806c
		x"2b6f0008", -- 18070
		x"fff6defc", -- 18074
		x"000c4efa", -- 18078
		x"001c2c5f", -- 1807c
		x"2b5ffff6", -- 18080
		x"7022b06d", -- 18084
		x"fffe6600", -- 18088
		x"00044e4a", -- 1808c
		x"3b7c0021", -- 18090
		x"fffe4e4a", -- 18094
		x"0cae0000", -- 18098
		x"0000fff8", -- 1809c
		x"6e00ff6e", -- 180a0
		x"2d7c0000", -- 180a4
		x"0100fff8", -- 180a8
		x"53aefff8", -- 180ac
		x"2f2dfff6", -- 180b0
		x"2f0e487a", -- 180b4
		x"001e2b4f", -- 180b8
		x"fff6206e", -- 180bc
		x"fff0116e", -- 180c0
		x"fffb003d", -- 180c4
		x"2b6f0008", -- 180c8
		x"fff6defc", -- 180cc
		x"000c4efa", -- 180d0
		x"00102c5f", -- 180d4
		x"2b5ffff6", -- 180d8
		x"3b7c0023", -- 180dc
		x"fffe4e4a", -- 180e0
		x"2f2dfff6", -- 180e4
		x"2f0e487a", -- 180e8
		x"002e2b4f", -- 180ec
		x"fff6206e", -- 180f0
		x"fff07000", -- 180f4
		x"1028003d", -- 180f8
		x"b0aefff8", -- 180fc
		x"6700000a", -- 18100
		x"3b7c0025", -- 18104
		x"fffe4e4a", -- 18108
		x"2b6f0008", -- 1810c
		x"fff6defc", -- 18110
		x"000c4efa", -- 18114
		x"001c2c5f", -- 18118
		x"2b5ffff6", -- 1811c
		x"7025b06d", -- 18120
		x"fffe6600", -- 18124
		x"00044e4a", -- 18128
		x"3b7c0024", -- 1812c
		x"fffe4e4a", -- 18130
		x"0cae0000", -- 18134
		x"0000fff8", -- 18138
		x"6e00ff6e", -- 1813c
		x"4a2e0008", -- 18140
		x"670000b6", -- 18144
		x"2d7c0000", -- 18148
		x"0100fff8", -- 1814c
		x"53aefff8", -- 18150
		x"598f2f2e", -- 18154
		x"fff82f3c", -- 18158
		x"00000030", -- 1815c
		x"4eb90000", -- 18160
		x"a9d44a9f", -- 18164
		x"66000086", -- 18168
		x"2f2dfff6", -- 1816c
		x"2f0e487a", -- 18170
		x"001e2b4f", -- 18174
		x"fff6206e", -- 18178
		x"fff0116e", -- 1817c
		x"fffb0005", -- 18180
		x"2b6f0008", -- 18184
		x"fff6defc", -- 18188
		x"000c4efa", -- 1818c
		x"00102c5f", -- 18190
		x"2b5ffff6", -- 18194
		x"3b7c0007", -- 18198
		x"fffe4e4a", -- 1819c
		x"2f2dfff6", -- 181a0
		x"2f0e487a", -- 181a4
		x"002e2b4f", -- 181a8
		x"fff6206e", -- 181ac
		x"fff07000", -- 181b0
		x"1028002b", -- 181b4
		x"b0aefff8", -- 181b8
		x"6700000a", -- 181bc
		x"3b7c0027", -- 181c0
		x"fffe4e4a", -- 181c4
		x"2b6f0008", -- 181c8
		x"fff6defc", -- 181cc
		x"000c4efa", -- 181d0
		x"001c2c5f", -- 181d4
		x"2b5ffff6", -- 181d8
		x"7027b06d", -- 181dc
		x"fffe6600", -- 181e0
		x"00044e4a", -- 181e4
		x"3b7c0026", -- 181e8
		x"fffe4e4a", -- 181ec
		x"0cae0000", -- 181f0
		x"0000fff8", -- 181f4
		x"6e00ff56", -- 181f8
		x"2f2dfff6", -- 181fc
		x"2f0e487a", -- 18200
		x"002a2b4f", -- 18204
		x"fff6206e", -- 18208
		x"fff07005", -- 1820c
		x"b028002d", -- 18210
		x"6700000a", -- 18214
		x"3b7c0029", -- 18218
		x"fffe4e4a", -- 1821c
		x"2b6f0008", -- 18220
		x"fff6defc", -- 18224
		x"000c4efa", -- 18228
		x"001c2c5f", -- 1822c
		x"2b5ffff6", -- 18230
		x"7029b06d", -- 18234
		x"fffe6600", -- 18238
		x"00044e4a", -- 1823c
		x"3b7c0028", -- 18240
		x"fffe4e4a", -- 18244
		x"2f2dfff6", -- 18248
		x"2f0e487a", -- 1824c
		x"001e2b4f", -- 18250
		x"fff6206e", -- 18254
		x"fff0117c", -- 18258
		x"ff01003d", -- 1825c
		x"2b6f0008", -- 18260
		x"fff6defc", -- 18264
		x"000c4efa", -- 18268
		x"00102c5f", -- 1826c
		x"2b5ffff6", -- 18270
		x"3b7c0023", -- 18274
		x"fffe4e4a", -- 18278
		x"2f2dfff6", -- 1827c
		x"2f0e487a", -- 18280
		x"002a2b4f", -- 18284
		x"fff6206e", -- 18288
		x"fff07001", -- 1828c
		x"b028002d", -- 18290
		x"6700000a", -- 18294
		x"3b7c0029", -- 18298
		x"fffe4e4a", -- 1829c
		x"2b6f0008", -- 182a0
		x"fff6defc", -- 182a4
		x"000c4efa", -- 182a8
		x"001c2c5f", -- 182ac
		x"2b5ffff6", -- 182b0
		x"7029b06d", -- 182b4
		x"fffe6600", -- 182b8
		x"00044e4a", -- 182bc
		x"3b7c0028", -- 182c0
		x"fffe4e4a", -- 182c4
		x"2f2dfff6", -- 182c8
		x"2f0e487a", -- 182cc
		x"001e2b4f", -- 182d0
		x"fff6206e", -- 182d4
		x"fff0117c", -- 182d8
		x"ff00003d", -- 182dc
		x"2b6f0008", -- 182e0
		x"fff6defc", -- 182e4
		x"000c4efa", -- 182e8
		x"00102c5f", -- 182ec
		x"2b5ffff6", -- 182f0
		x"3b7c0023", -- 182f4
		x"fffe4e4a", -- 182f8
		x"2f2dfff6", -- 182fc
		x"2f0e487a", -- 18300
		x"001e2b4f", -- 18304
		x"fff6206e", -- 18308
		x"fff0117c", -- 1830c
		x"ffff0029", -- 18310
		x"2b6f0008", -- 18314
		x"fff6defc", -- 18318
		x"000c4efa", -- 1831c
		x"00102c5f", -- 18320
		x"2b5ffff6", -- 18324
		x"3b7c002a", -- 18328
		x"fffe4e4a", -- 1832c
		x"2f2dfff6", -- 18330
		x"2f0e487a", -- 18334
		x"00282b4f", -- 18338
		x"fff6206e", -- 1833c
		x"fff04a28", -- 18340
		x"00296700", -- 18344
		x"000a3b7c", -- 18348
		x"002cfffe", -- 1834c
		x"4e4a2b6f", -- 18350
		x"0008fff6", -- 18354
		x"defc000c", -- 18358
		x"4efa001c", -- 1835c
		x"2c5f2b5f", -- 18360
		x"fff6702c", -- 18364
		x"b06dfffe", -- 18368
		x"66000004", -- 1836c
		x"4e4a3b7c", -- 18370
		x"002bfffe", -- 18374
		x"4e4a2f2d", -- 18378
		x"fff62f0e", -- 1837c
		x"487a0028", -- 18380
		x"2b4ffff6", -- 18384
		x"206efff0", -- 18388
		x"4a28002f", -- 1838c
		x"6700000a", -- 18390
		x"3b7c002e", -- 18394
		x"fffe4e4a", -- 18398
		x"2b6f0008", -- 1839c
		x"fff6defc", -- 183a0
		x"000c4efa", -- 183a4
		x"001c2c5f", -- 183a8
		x"2b5ffff6", -- 183ac
		x"702eb06d", -- 183b0
		x"fffe6600", -- 183b4
		x"00044e4a", -- 183b8
		x"3b7c002d", -- 183bc
		x"fffe4e4a", -- 183c0
		x"2f2dfff6", -- 183c4
		x"2f0e487a", -- 183c8
		x"00282b4f", -- 183cc
		x"fff6206e", -- 183d0
		x"fff04a28", -- 183d4
		x"00336700", -- 183d8
		x"000a3b7c", -- 183dc
		x"0030fffe", -- 183e0
		x"4e4a2b6f", -- 183e4
		x"0008fff6", -- 183e8
		x"defc000c", -- 183ec
		x"4efa001c", -- 183f0
		x"2c5f2b5f", -- 183f4
		x"fff67030", -- 183f8
		x"b06dfffe", -- 183fc
		x"66000004", -- 18400
		x"4e4a3b7c", -- 18404
		x"002ffffe", -- 18408
		x"4e4a2f0e", -- 1840c
		x"4ebaf732", -- 18410
		x"4e5e205f", -- 18414
		x"5c4f4ed0", -- 18418
		x"4e750000", -- 1841c
		x"4e56fff2", -- 18420
		x"2f2e0008", -- 18424
		x"42274eb9", -- 18428
		x"00016788", -- 1842c
		x"2d6e0008", -- 18430
		x"fff22f2d", -- 18434
		x"fff62f0e", -- 18438
		x"487a0100", -- 1843c
		x"2b4ffff6", -- 18440
		x"206efff2", -- 18444
		x"117cff00", -- 18448
		x"00232d7c", -- 1844c
		x"ffffffff", -- 18450
		x"fff852ae", -- 18454
		x"fff8206e", -- 18458
		x"fff2117c", -- 1845c
		x"ff01003b", -- 18460
		x"117cff04", -- 18464
		x"003d116e", -- 18468
		x"fffb0037", -- 1846c
		x"117cff20", -- 18470
		x"00252d7c", -- 18474
		x"00000080", -- 18478
		x"fffc4aae", -- 1847c
		x"fffc6f00", -- 18480
		x"005e202e", -- 18484
		x"fffc0280", -- 18488
		x"0000000f", -- 1848c
		x"4a806600", -- 18490
		x"0048206e", -- 18494
		x"fff27000", -- 18498
		x"10280029", -- 1849c
		x"3d40fff6", -- 184a0
		x"598f302e", -- 184a4
		x"fff648c0", -- 184a8
		x"2f00598f", -- 184ac
		x"2f3c0000", -- 184b0
		x"00044eb9", -- 184b4
		x"0000a9de", -- 184b8
		x"4eb90000", -- 184bc
		x"a9d44a9f", -- 184c0
		x"6700000a", -- 184c4
		x"3b7c002c", -- 184c8
		x"fffe4e4a", -- 184cc
		x"4a6efff6", -- 184d0
		x"67000006", -- 184d4
		x"42aefffc", -- 184d8
		x"53aefffc", -- 184dc
		x"609c4aae", -- 184e0
		x"fffc6c00", -- 184e4
		x"002a206e", -- 184e8
		x"fff27000", -- 184ec
		x"10280005", -- 184f0
		x"3d40fff6", -- 184f4
		x"302efff6", -- 184f8
		x"48c0b0ae", -- 184fc
		x"fff86700", -- 18500
		x"000a3b7c", -- 18504
		x"001cfffe", -- 18508
		x"4e4a6000", -- 1850c
		x"000a3b7c", -- 18510
		x"0033fffe", -- 18514
		x"4e4a0cae", -- 18518
		x"000000ff", -- 1851c
		x"fff86d00", -- 18520
		x"ff32206e", -- 18524
		x"fff2117c", -- 18528
		x"ff800023", -- 1852c
		x"2b6f0008", -- 18530
		x"fff6defc", -- 18534
		x"000c4efa", -- 18538
		x"00342c5f", -- 1853c
		x"2b5ffff6", -- 18540
		x"206efff2", -- 18544
		x"117cff80", -- 18548
		x"0023302d", -- 1854c
		x"fffe48c0", -- 18550
		x"2f00487a", -- 18554
		x"001e4eb9", -- 18558
		x"000081b4", -- 1855c
		x"4a1f6700", -- 18560
		x"00044e4a", -- 18564
		x"3b7c0032", -- 18568
		x"fffe4e4a", -- 1856c
		x"4e5e2e9f", -- 18570
		x"4e750008", -- 18574
		x"00000008", -- 18578
		x"00081000", -- 1857c
		x"00004e56", -- 18580
		x"fff62f2e", -- 18584
		x"000c4227", -- 18588
		x"4eb90001", -- 1858c
		x"67883d7c", -- 18590
		x"0011fffe", -- 18594
		x"4a2e000a", -- 18598
		x"67000008", -- 1859c
		x"066e0020", -- 185a0
		x"fffe2d6e", -- 185a4
		x"000cfff6", -- 185a8
		x"2f2dfff6", -- 185ac
		x"2f0e487a", -- 185b0
		x"002a2b4f", -- 185b4
		x"fff6302e", -- 185b8
		x"fffed07c", -- 185bc
		x"0080206e", -- 185c0
		x"fff61140", -- 185c4
		x"0023116e", -- 185c8
		x"ffff0023", -- 185cc
		x"2b6f0008", -- 185d0
		x"fff6defc", -- 185d4
		x"000c4efa", -- 185d8
		x"00102c5f", -- 185dc
		x"2b5ffff6", -- 185e0
		x"3b7c000e", -- 185e4
		x"fffe4e4a", -- 185e8
		x"4a2e000a", -- 185ec
		x"67000014", -- 185f0
		x"2d6e000c", -- 185f4
		x"fffa06ae", -- 185f8
		x"0000002a", -- 185fc
		x"fffa6000", -- 18600
		x"000c2d6e", -- 18604
		x"000cfffa", -- 18608
		x"58aefffa", -- 1860c
		x"558f2f2e", -- 18610
		x"000c2f2e", -- 18614
		x"fffa3f2e", -- 18618
		x"00084eb9", -- 1861c
		x"00016e9a", -- 18620
		x"4a1f6700", -- 18624
		x"002c2f2e", -- 18628
		x"000c2f2e", -- 1862c
		x"fffa4eb9", -- 18630
		x"00017004", -- 18634
		x"2f2e000c", -- 18638
		x"2f2efffa", -- 1863c
		x"4eb90001", -- 18640
		x"714c2f2e", -- 18644
		x"000c2f2e", -- 18648
		x"fffa4eb9", -- 1864c
		x"000176d6", -- 18650
		x"4e5e205f", -- 18654
		x"504f4ed0", -- 18658
		x"00004e56", -- 1865c
		x"ffec2d6e", -- 18660
		x"000cfff4", -- 18664
		x"206efff4", -- 18668
		x"2d680004", -- 1866c
		x"fff02d68", -- 18670
		x"0018ffec", -- 18674
		x"2d680004", -- 18678
		x"fffc58ae", -- 1867c
		x"fffc2f28", -- 18680
		x"00044227", -- 18684
		x"4eb90001", -- 18688
		x"67882f2d", -- 1868c
		x"fff62f0e", -- 18690
		x"487a0024", -- 18694
		x"2b4ffff6", -- 18698
		x"206efff0", -- 1869c
		x"117cff91", -- 186a0
		x"0023117c", -- 186a4
		x"ff110023", -- 186a8
		x"2b6f0008", -- 186ac
		x"fff6defc", -- 186b0
		x"000c4efa", -- 186b4
		x"00102c5f", -- 186b8
		x"2b5ffff6", -- 186bc
		x"3b7c000e", -- 186c0
		x"fffe4e4a", -- 186c4
		x"558f206e", -- 186c8
		x"fff42f28", -- 186cc
		x"00042f2e", -- 186d0
		x"fffc3f2e", -- 186d4
		x"00084eb9", -- 186d8
		x"00016e9a", -- 186dc
		x"4a1f6700", -- 186e0
		x"004a2d7c", -- 186e4
		x"ffffffff", -- 186e8
		x"fff852ae", -- 186ec
		x"fff8206e", -- 186f0
		x"fff42f28", -- 186f4
		x"0004226e", -- 186f8
		x"ffec2f29", -- 186fc
		x"00021f2e", -- 18700
		x"000a4227", -- 18704
		x"2f2efff8", -- 18708
		x"4eb90001", -- 1870c
		x"74de0cae", -- 18710
		x"00000001", -- 18714
		x"fff86dd2", -- 18718
		x"206efff4", -- 1871c
		x"2f280004", -- 18720
		x"2f2efffc", -- 18724
		x"4eb90001", -- 18728
		x"76d64e5e", -- 1872c
		x"205f504f", -- 18730
		x"4ed04e75", -- 18734
		x"00000000", -- 18738
		x"00080000", -- 1873c
		x"00090000", -- 18740
		x"01050e0c", -- 18744
		x"00000000", -- 18748
		x"00000000", -- 1874c
		x"00000000", -- 18750
		x"00000102", -- 18754
		x"4dfa0068", -- 18758
		x"41f90040", -- 1875c
		x"8000ba28", -- 18760
		x"0001662a", -- 18764
		x"12280003", -- 18768
		x"020100f0", -- 1876c
		x"0c010010", -- 18770
		x"661c48e7", -- 18774
		x"ee804284", -- 18778
		x"09080005", -- 1877c
		x"e38c4eb9", -- 18780
		x"00004eaa", -- 18784
		x"4cdf0177", -- 18788
		x"4a43661a", -- 1878c
		x"60360c28", -- 18790
		x"00ff0001", -- 18794
		x"67284281", -- 18798
		x"03080005", -- 1879c
		x"e3896706", -- 187a0
		x"41f01800", -- 187a4
		x"60b808f8", -- 187a8
		x"0000fed9", -- 187ac
		x"0c050001", -- 187b0
		x"66044287", -- 187b4
		x"60080c05", -- 187b8
		x"00036602", -- 187bc
		x"4286023c", -- 187c0
		x"001b4e75", -- 187c4
		x"003c0004", -- 187c8
		x"4e751228", -- 187cc
		x"000067ee", -- 187d0
		x"0c010001", -- 187d4
		x"6606b028", -- 187d8
		x"000867e8", -- 187dc
		x"42811228", -- 187e0
		x"0002e349", -- 187e4
		x"67c041f0", -- 187e8
		x"100060de", -- 187ec
		x"2878fed4", -- 187f0
		x"0200007f", -- 187f4
		x"14000202", -- 187f8
		x"001f4a28", -- 187fc
		x"000067be", -- 18800
		x"0c280001", -- 18804
		x"00006618", -- 18808
		x"b0280010", -- 1880c
		x"67b61628", -- 18810
		x"00100203", -- 18814
		x"001fb403", -- 18818
		x"67aab028", -- 1881c
		x"000e67a4", -- 18820
		x"42411228", -- 18824
		x"0002e349", -- 18828
		x"6700ff7c", -- 1882c
		x"41f01000", -- 18830
		x"60c84a29", -- 18834
		x"00006786", -- 18838
		x"01490006", -- 1883c
		x"b2806784", -- 18840
		x"42801029", -- 18844
		x"0002e348", -- 18848
		x"6700ff5c", -- 1884c
		x"41f10000", -- 18850
		x"60e04dfa", -- 18854
		x"00c04280", -- 18858
		x"10280004", -- 1885c
		x"e34841f0", -- 18860
		x"00ff4282", -- 18864
		x"42832441", -- 18868
		x"36184a03", -- 1886c
		x"670000a6", -- 18870
		x"0c030001", -- 18874
		x"66083418", -- 18878
		x"024200ff", -- 1887c
		x"60ea0c03", -- 18880
		x"00026608", -- 18884
		x"05080001", -- 18888
		x"584860dc", -- 1888c
		x"0c030003", -- 18890
		x"66083818", -- 18894
		x"15842800", -- 18898
		x"60ce0c03", -- 1889c
		x"0004661c", -- 188a0
		x"38180244", -- 188a4
		x"00ff45f2", -- 188a8
		x"28006008", -- 188ac
		x"14a80001", -- 188b0
		x"5448544a", -- 188b4
		x"51ccfff6", -- 188b8
		x"244160ac", -- 188bc
		x"0c030005", -- 188c0
		x"661a3818", -- 188c4
		x"024400ff", -- 188c8
		x"45f22800", -- 188cc
		x"30186004", -- 188d0
		x"1480544a", -- 188d4
		x"51ccfffa", -- 188d8
		x"2441608c", -- 188dc
		x"0c030006", -- 188e0
		x"66044a11", -- 188e4
		x"60820c03", -- 188e8
		x"00076606", -- 188ec
		x"12916000", -- 188f0
		x"ff780c03", -- 188f4
		x"0008660a", -- 188f8
		x"38188932", -- 188fc
		x"28006000", -- 18900
		x"ff680c03", -- 18904
		x"00096600", -- 18908
		x"fe9e3818", -- 1890c
		x"c9322800", -- 18910
		x"6000ff56", -- 18914
		x"4e754dfa", -- 18918
		x"003a41f9", -- 1891c
		x"00400011", -- 18920
		x"42801010", -- 18924
		x"0c000060", -- 18928
		x"6d284840", -- 1892c
		x"22401229", -- 18930
		x"00010201", -- 18934
		x"007f0c01", -- 18938
		x"00156616", -- 1893c
		x"d3fc0000", -- 18940
		x"c00145fa", -- 18944
		x"fdf0741f", -- 18948
		x"129a43e9", -- 1894c
		x"000251ca", -- 18950
		x"fff841e8", -- 18954
		x"0002b1fc", -- 18958
		x"00400041", -- 1895c
		x"66c24dfa", -- 18960
		x"01b80839", -- 18964
		x"00030040", -- 18968
		x"00036700", -- 1896c
		x"01ac4287", -- 18970
		x"7a016100", -- 18974
		x"fde06670", -- 18978
		x"2e084dfa", -- 1897c
		x"000c43f9", -- 18980
		x"00400011", -- 18984
		x"10111280", -- 18988
		x"43e90002", -- 1898c
		x"b3fc0040", -- 18990
		x"004166f0", -- 18994
		x"4dfa0024", -- 18998
		x"41e80015", -- 1899c
		x"43f90040", -- 189a0
		x"00101028", -- 189a4
		x"0000672a", -- 189a8
		x"0c000001", -- 189ac
		x"660c4281", -- 189b0
		x"12280012", -- 189b4
		x"13a80008", -- 189b8
		x"10004281", -- 189bc
		x"12280002", -- 189c0
		x"e3496706", -- 189c4
		x"41f01000", -- 189c8
		x"60d808f8", -- 189cc
		x"0000fed9", -- 189d0
		x"42874dfa", -- 189d4
		x"000a43f9", -- 189d8
		x"00400011", -- 189dc
		x"10115449", -- 189e0
		x"b3fc0040", -- 189e4
		x"004166f4", -- 189e8
		x"42861a3c", -- 189ec
		x"00036100", -- 189f0
		x"fd646602", -- 189f4
		x"2c084dfa", -- 189f8
		x"009243f9", -- 189fc
		x"00400011", -- 18a00
		x"10114a87", -- 18a04
		x"673e2047", -- 18a08
		x"7a0141e8", -- 18a0c
		x"00156100", -- 18a10
		x"fdba6630", -- 18a14
		x"0c000060", -- 18a18
		x"6d5c0348", -- 18a1c
		x"00062441", -- 18a20
		x"102a0001", -- 18a24
		x"0200007f", -- 18a28
		x"b0280010", -- 18a2c
		x"6748b028", -- 18a30
		x"000e6742", -- 18a34
		x"0200001f", -- 18a38
		x"1228000e", -- 18a3c
		x"0201001f", -- 18a40
		x"b0016732", -- 18a44
		x"4a866700", -- 18a48
		x"00422046", -- 18a4c
		x"7a0341e8", -- 18a50
		x"00150c00", -- 18a54
		x"00606d16", -- 18a58
		x"42811200", -- 18a5c
		x"48412441", -- 18a60
		x"102a0001", -- 18a64
		x"6100fd86", -- 18a68
		x"670c6000", -- 18a6c
		x"001e6100", -- 18a70
		x"fd5a6600", -- 18a74
		x"00160348", -- 18a78
		x"00064a81", -- 18a7c
		x"66041211", -- 18a80
		x"48411291", -- 18a84
		x"6100fdcc", -- 18a88
		x"4a114dfa", -- 18a8c
		x"fffe5449", -- 18a90
		x"b3fc0040", -- 18a94
		x"00416600", -- 18a98
		x"ff684238", -- 18a9c
		x"fdcc4a87", -- 18aa0
		x"67482047", -- 18aa4
		x"7a0141e8", -- 18aa8
		x"00154a28", -- 18aac
		x"0000673a", -- 18ab0
		x"0c100002", -- 18ab4
		x"66240348", -- 18ab8
		x"00064a38", -- 18abc
		x"fdcc6712", -- 18ac0
		x"4a87670e", -- 18ac4
		x"22477a01", -- 18ac8
		x"43e90015", -- 18acc
		x"6100fd64", -- 18ad0
		x"67082248", -- 18ad4
		x"6100fd7c", -- 18ad8
		x"20494280", -- 18adc
		x"10280002", -- 18ae0
		x"e348671e", -- 18ae4
		x"41f00000", -- 18ae8
		x"60c04a38", -- 18aec
		x"fdcc661e", -- 18af0
		x"4638fdcc", -- 18af4
		x"4a866716", -- 18af8
		x"20467a03", -- 18afc
		x"41e80015", -- 18b00
		x"60a808f8", -- 18b04
		x"0000fed9", -- 18b08
		x"4a38fdcc", -- 18b0c
		x"67dc2878", -- 18b10
		x"fed408ec", -- 18b14
		x"0004000a", -- 18b18
		x"4e750001", -- 18b1c
		x"8b3a0001", -- 18b20
		x"00018c6c", -- 18b24
		x"00000000", -- 18b28
		x"00000000", -- 18b2c
		x"00000000", -- 18b30
		x"20202050", -- 18b34
		x"00000001", -- 18b38
		x"8b560001", -- 18b3c
		x"0001926c", -- 18b40
		x"00000000", -- 18b44
		x"00000000", -- 18b48
		x"00000000", -- 18b4c
		x"20202054", -- 18b50
		x"00000001", -- 18b54
		x"8b720001", -- 18b58
		x"00018f7a", -- 18b5c
		x"00000000", -- 18b60
		x"00000000", -- 18b64
		x"00000000", -- 18b68
		x"2020204c", -- 18b6c
		x"00000001", -- 18b70
		x"8b8e0001", -- 18b74
		x"0001be16", -- 18b78
		x"00000000", -- 18b7c
		x"00000000", -- 18b80
		x"00000000", -- 18b84
		x"20202043", -- 18b88
		x"00000001", -- 18b8c
		x"8baa0001", -- 18b90
		x"00018c74", -- 18b94
		x"00000000", -- 18b98
		x"00000000", -- 18b9c
		x"00000000", -- 18ba0
		x"20202020", -- 18ba4
		x"00000000", -- 18ba8
		x"00000001", -- 18bac
		x"00018c98", -- 18bb0
		x"00000000", -- 18bb4
		x"00000000", -- 18bb8
		x"00000000", -- 18bbc
		x"20202020", -- 18bc0
		x"000048e7", -- 18bc4
		x"fffe2878", -- 18bc8
		x"fed44eb9", -- 18bcc
		x"00006d78", -- 18bd0
		x"4a2c00c0", -- 18bd4
		x"6d00008c", -- 18bd8
		x"202c00ca", -- 18bdc
		x"08ac0001", -- 18be0
		x"00c06606", -- 18be4
		x"103c0020", -- 18be8
		x"e0980c00", -- 18bec
		x"0020660a", -- 18bf0
		x"e0980c00", -- 18bf4
		x"00206602", -- 18bf8
		x"e098206c", -- 18bfc
		x"00c6082c", -- 18c00
		x"0002000b", -- 18c04
		x"671e11c0", -- 18c08
		x"fdd2197c", -- 18c0c
		x"000300ba", -- 18c10
		x"08ec0000", -- 18c14
		x"00c008ec", -- 18c18
		x"000200c0", -- 18c1c
		x"08ac0002", -- 18c20
		x"000b601a", -- 18c24
		x"122c00c1", -- 18c28
		x"c2280004", -- 18c2c
		x"b2280004", -- 18c30
		x"6626b0a8", -- 18c34
		x"00166620", -- 18c38
		x"22680006", -- 18c3c
		x"4e912878", -- 18c40
		x"fed4197c", -- 18c44
		x"000300bb", -- 18c48
		x"08ec0003", -- 18c4c
		x"00c008ec", -- 18c50
		x"000700c0", -- 18c54
		x"6000ff74", -- 18c58
		x"22280000", -- 18c5c
		x"67da2041", -- 18c60
		x"60c24cdf", -- 18c64
		x"7fff4e75", -- 18c68
		x"08ec0002", -- 18c6c
		x"005c4e75", -- 18c70
		x"08ac0002", -- 18c74
		x"005c661a", -- 18c78
		x"08ec0007", -- 18c7c
		x"000a397c", -- 18c80
		x"0020032c", -- 18c84
		x"082c0006", -- 18c88
		x"000a6606", -- 18c8c
		x"4eb90000", -- 18c90
		x"58304e75", -- 18c94
		x"b03c0041", -- 18c98
		x"6570b03c", -- 18c9c
		x"005a630c", -- 18ca0
		x"b03c0061", -- 18ca4
		x"6564b03c", -- 18ca8
		x"007a625e", -- 18cac
		x"1600e098", -- 18cb0
		x"b03c0030", -- 18cb4
		x"65000054", -- 18cb8
		x"b03c0039", -- 18cbc
		x"6200004c", -- 18cc0
		x"42811200", -- 18cc4
		x"04410030", -- 18cc8
		x"e0980c00", -- 18ccc
		x"0020671e", -- 18cd0
		x"b03c0030", -- 18cd4
		x"65000034", -- 18cd8
		x"b03c0039", -- 18cdc
		x"6200002c", -- 18ce0
		x"42821400", -- 18ce4
		x"04420030", -- 18ce8
		x"c4fc000a", -- 18cec
		x"d2821941", -- 18cf0
		x"032c1943", -- 18cf4
		x"032d08ec", -- 18cf8
		x"0007000a", -- 18cfc
		x"082c0006", -- 18d00
		x"000a6606", -- 18d04
		x"4eb90000", -- 18d08
		x"58304e75", -- 18d0c
		x"205f225f", -- 18d10
		x"245f265f", -- 18d14
		x"2f082878", -- 18d18
		x"fed4206c", -- 18d1c
		x"00b62010", -- 18d20
		x"0c802020", -- 18d24
		x"2020671a", -- 18d28
		x"0c802020", -- 18d2c
		x"20596708", -- 18d30
		x"0c802020", -- 18d34
		x"204e660e", -- 18d38
		x"266dfff0", -- 18d3c
		x"4e9312bc", -- 18d40
		x"000114bc", -- 18d44
		x"00014e75", -- 18d48
		x"00018d84", -- 18d4c
		x"00005479", -- 18d50
		x"70652059", -- 18d54
		x"206f7220", -- 18d58
		x"4e20454e", -- 18d5c
		x"54455220", -- 18d60
		x"3f200000", -- 18d64
		x"00018d84", -- 18d68
		x"00005479", -- 18d6c
		x"70652059", -- 18d70
		x"206f7220", -- 18d74
		x"4e205245", -- 18d78
		x"5455524e", -- 18d7c
		x"203f2000", -- 18d80
		x"00018d8c", -- 18d84
		x"00032000", -- 18d88
		x"00000000", -- 18d8c
		x"00010001", -- 18d90
		x"8d100000", -- 18d94
		x"00000000", -- 18d98
		x"00000000", -- 18d9c
		x"00002020", -- 18da0
		x"2020ff63", -- 18da4
		x"205f225f", -- 18da8
		x"245f265f", -- 18dac
		x"2f084a11", -- 18db0
		x"672441eb", -- 18db4
		x"001a3010", -- 18db8
		x"6c0441f5", -- 18dbc
		x"0000226b", -- 18dc0
		x"000e10d9", -- 18dc4
		x"66fc5388", -- 18dc8
		x"266b0012", -- 18dcc
		x"42804e93", -- 18dd0
		x"10c04210", -- 18dd4
		x"4e752f09", -- 18dd8
		x"41edff63", -- 18ddc
		x"43eb001a", -- 18de0
		x"30116e04", -- 18de4
		x"43f50000", -- 18de8
		x"10d966fc", -- 18dec
		x"2b6b0012", -- 18df0
		x"fff0225f", -- 18df4
		x"41faff6e", -- 18df8
		x"4a2c00a9", -- 18dfc
		x"660441fa", -- 18e00
		x"ff482f08", -- 18e04
		x"422712bc", -- 18e08
		x"00012f09", -- 18e0c
		x"4eba06ae", -- 18e10
		x"4e752278", -- 18e14
		x"fed40829", -- 18e18
		x"0004000b", -- 18e1c
		x"671e007c", -- 18e20
		x"070049f8", -- 18e24
		x"f738204c", -- 18e28
		x"45f8fac0", -- 18e2c
		x"20d9b5c8", -- 18e30
		x"62fa21cc", -- 18e34
		x"fed408ac", -- 18e38
		x"0004000b", -- 18e3c
		x"4ef90000", -- 18e40
		x"074e205f", -- 18e44
		x"225f245f", -- 18e48
		x"245f12bc", -- 18e4c
		x"00012878", -- 18e50
		x"fed408b8", -- 18e54
		x"0006fed2", -- 18e58
		x"08ac0000", -- 18e5c
		x"000a08ec", -- 18e60
		x"0001000b", -- 18e64
		x"08ac0000", -- 18e68
		x"000b4ed0", -- 18e6c
		x"205f225f", -- 18e70
		x"245f265f", -- 18e74
		x"2f082878", -- 18e78
		x"fed4206c", -- 18e7c
		x"00b62010", -- 18e80
		x"0c802020", -- 18e84
		x"2020671a", -- 18e88
		x"0c802020", -- 18e8c
		x"35306708", -- 18e90
		x"0c802020", -- 18e94
		x"3630660e", -- 18e98
		x"266dfff0", -- 18e9c
		x"4e9312bc", -- 18ea0
		x"000114bc", -- 18ea4
		x"00014e75", -- 18ea8
		x"00018ee8", -- 18eac
		x"00005479", -- 18eb0
		x"70652035", -- 18eb4
		x"30206f72", -- 18eb8
		x"20363020", -- 18ebc
		x"454e5445", -- 18ec0
		x"52203f20", -- 18ec4
		x"00000001", -- 18ec8
		x"8ee80000", -- 18ecc
		x"54797065", -- 18ed0
		x"20353020", -- 18ed4
		x"6f722036", -- 18ed8
		x"30205245", -- 18edc
		x"5455524e", -- 18ee0
		x"203f2000", -- 18ee4
		x"00018ef0", -- 18ee8
		x"00032000", -- 18eec
		x"00000000", -- 18ef0
		x"00010001", -- 18ef4
		x"8e700000", -- 18ef8
		x"00000000", -- 18efc
		x"00000000", -- 18f00
		x"00002020", -- 18f04
		x"2020ff63", -- 18f08
		x"205f225f", -- 18f0c
		x"245f265f", -- 18f10
		x"2f084a11", -- 18f14
		x"672441eb", -- 18f18
		x"001a3010", -- 18f1c
		x"6c0441f5", -- 18f20
		x"0000226b", -- 18f24
		x"000e10d9", -- 18f28
		x"66fc5388", -- 18f2c
		x"266b0012", -- 18f30
		x"42804e93", -- 18f34
		x"30c04210", -- 18f38
		x"4e752f09", -- 18f3c
		x"41edff63", -- 18f40
		x"43eb001a", -- 18f44
		x"30116e04", -- 18f48
		x"43f50000", -- 18f4c
		x"10d966fc", -- 18f50
		x"2b6b0012", -- 18f54
		x"fff0225f", -- 18f58
		x"41faff6c", -- 18f5c
		x"4a2c00a9", -- 18f60
		x"660441fa", -- 18f64
		x"ff442f08", -- 18f68
		x"422712bc", -- 18f6c
		x"00012f09", -- 18f70
		x"4eba054a", -- 18f74
		x"4e75082c", -- 18f78
		x"0001005c", -- 18f7c
		x"67164a2c", -- 18f80
		x"005d66f0", -- 18f84
		x"197c0001", -- 18f88
		x"005d297c", -- 18f8c
		x"00018f98", -- 18f90
		x"00c260e0", -- 18f94
		x"08f80001", -- 18f98
		x"fed94efa", -- 18f9c
		x"fe760001", -- 18fa0
		x"8fd80000", -- 18fa4
		x"54797065", -- 18fa8
		x"205b6b65", -- 18fac
		x"795d2045", -- 18fb0
		x"4e544552", -- 18fb4
		x"203f2000", -- 18fb8
		x"00018fd8", -- 18fbc
		x"00005479", -- 18fc0
		x"7065205b", -- 18fc4
		x"6b65795d", -- 18fc8
		x"20524554", -- 18fcc
		x"55524e20", -- 18fd0
		x"3f200000", -- 18fd4
		x"00018ff6", -- 18fd8
		x"00032020", -- 18fdc
		x"20205365", -- 18fe0
		x"6c662054", -- 18fe4
		x"65737420", -- 18fe8
		x"436f6e74", -- 18fec
		x"726f6c73", -- 18ff0
		x"00000001", -- 18ff4
		x"90180003", -- 18ff8
		x"4b657973", -- 18ffc
		x"20546573", -- 19000
		x"74204f70", -- 19004
		x"74696f6e", -- 19008
		x"20202053", -- 1900c
		x"656c6563", -- 19010
		x"74656400", -- 19014
		x"0001907a", -- 19018
		x"00032d2d", -- 1901c
		x"2d2d2d2d", -- 19020
		x"2d2d2d2d", -- 19024
		x"2d2d2d2d", -- 19028
		x"2d2d2d2d", -- 1902c
		x"2d2d2d2d", -- 19030
		x"2d2d2d2d", -- 19034
		x"2d002020", -- 19038
		x"31202043", -- 1903c
		x"6f6e7469", -- 19040
		x"6e756f75", -- 19044
		x"73202020", -- 19048
		x"20202020", -- 1904c
		x"20202000", -- 19050
		x"4a00660e", -- 19054
		x"70590838", -- 19058
		x"0006fed2", -- 1905c
		x"6602704e", -- 19060
		x"4e7508b8", -- 19064
		x"0006fed2", -- 19068
		x"0c00004e", -- 1906c
		x"67f208f8", -- 19070
		x"0006fed2", -- 19074
		x"4e750001", -- 19078
		x"90de0002", -- 1907c
		x"00018da8", -- 19080
		x"00000000", -- 19084
		x"0001903a", -- 19088
		x"00019054", -- 1908c
		x"20202031", -- 19090
		x"ffd32020", -- 19094
		x"32202045", -- 19098
		x"7874656e", -- 1909c
		x"64656420", -- 190a0
		x"20202020", -- 190a4
		x"20202020", -- 190a8
		x"20202000", -- 190ac
		x"2f0c2878", -- 190b0
		x"fed44a00", -- 190b4
		x"66107059", -- 190b8
		x"082c0000", -- 190bc
		x"000a6602", -- 190c0
		x"704e285f", -- 190c4
		x"4e7508ac", -- 190c8
		x"0000000a", -- 190cc
		x"0c00004e", -- 190d0
		x"67f008ec", -- 190d4
		x"0000000a", -- 190d8
		x"60e80001", -- 190dc
		x"91420002", -- 190e0
		x"00018da8", -- 190e4
		x"00000000", -- 190e8
		x"00019096", -- 190ec
		x"000190b0", -- 190f0
		x"20202032", -- 190f4
		x"ffb72020", -- 190f8
		x"33202054", -- 190fc
		x"65737420", -- 19100
		x"4d656d6f", -- 19104
		x"72792020", -- 19108
		x"20202020", -- 1910c
		x"20202000", -- 19110
		x"2f0c2878", -- 19114
		x"fed44a00", -- 19118
		x"66107059", -- 1911c
		x"082c0001", -- 19120
		x"000b6602", -- 19124
		x"704e285f", -- 19128
		x"4e7508ac", -- 1912c
		x"0001000b", -- 19130
		x"0c00004e", -- 19134
		x"67f008ec", -- 19138
		x"0001000b", -- 1913c
		x"60e80001", -- 19140
		x"91aa0002", -- 19144
		x"00018da8", -- 19148
		x"00000000", -- 1914c
		x"000190fa", -- 19150
		x"00019114", -- 19154
		x"20202033", -- 19158
		x"ff9b2020", -- 1915c
		x"34202035", -- 19160
		x"302f3630", -- 19164
		x"20487a20", -- 19168
		x"43525420", -- 1916c
		x"20202020", -- 19170
		x"20200000", -- 19174
		x"2f0c2878", -- 19178
		x"fed44a00", -- 1917c
		x"6614303c", -- 19180
		x"3530082c", -- 19184
		x"0000000b", -- 19188
		x"6604303c", -- 1918c
		x"3630285f", -- 19190
		x"4e7508ac", -- 19194
		x"0000000b", -- 19198
		x"0c403630", -- 1919c
		x"67f008ec", -- 191a0
		x"0000000b", -- 191a4
		x"60e80001", -- 191a8
		x"91c60102", -- 191ac
		x"00018f0c", -- 191b0
		x"00000000", -- 191b4
		x"0001915e", -- 191b8
		x"00019178", -- 191bc
		x"20202034", -- 191c0
		x"ff7f0001", -- 191c4
		x"91ce0003", -- 191c8
		x"20000001", -- 191cc
		x"91fa0001", -- 191d0
		x"00018e46", -- 191d4
		x"00000000", -- 191d8
		x"00000000", -- 191dc
		x"00000000", -- 191e0
		x"20202044", -- 191e4
		x"20204420", -- 191e8
		x"20736574", -- 191ec
		x"20446566", -- 191f0
		x"61756c74", -- 191f4
		x"73000001", -- 191f8
		x"92240001", -- 191fc
		x"00018e16", -- 19200
		x"00000000", -- 19204
		x"00000000", -- 19208
		x"00000000", -- 1920c
		x"20202052", -- 19210
		x"20205220", -- 19214
		x"2052756e", -- 19218
		x"20746573", -- 1921c
		x"74730000", -- 19220
		x"00000000", -- 19224
		x"00010001", -- 19228
		x"8c960000", -- 1922c
		x"00000000", -- 19230
		x"00000000", -- 19234
		x"00002020", -- 19238
		x"20202d2d", -- 1923c
		x"2d2d2d2d", -- 19240
		x"2d2d2d2d", -- 19244
		x"2d2d2d2d", -- 19248
		x"2d2d2d2d", -- 1924c
		x"2d2d2d2d", -- 19250
		x"2d2d2d2d", -- 19254
		x"2d002f0c", -- 19258
		x"2878fed4", -- 1925c
		x"082c0001", -- 19260
		x"005c6726", -- 19264
		x"285f4e75", -- 19268
		x"082c0001", -- 1926c
		x"005c671a", -- 19270
		x"4a2c005d", -- 19274
		x"660000be", -- 19278
		x"197c0001", -- 1927c
		x"005d297c", -- 19280
		x"0001925a", -- 19284
		x"00c26000", -- 19288
		x"00ac007c", -- 1928c
		x"07004ff8", -- 19290
		x"fdac2878", -- 19294
		x"fed4297c", -- 19298
		x"00018c96", -- 1929c
		x"00c241ec", -- 192a0
		x"00ca2948", -- 192a4
		x"00b6422c", -- 192a8
		x"00c0197c", -- 192ac
		x"000300ba", -- 192b0
		x"08ec0000", -- 192b4
		x"00c008ec", -- 192b8
		x"000200c0", -- 192bc
		x"08d40004", -- 192c0
		x"08ec0007", -- 192c4
		x"00c04eb9", -- 192c8
		x"00006d78", -- 192cc
		x"027cf0ff", -- 192d0
		x"082c0004", -- 192d4
		x"000b6606", -- 192d8
		x"294c0330", -- 192dc
		x"6008297c", -- 192e0
		x"fffffac0", -- 192e4
		x"03302a6c", -- 192e8
		x"033006ac", -- 192ec
		x"ffffff63", -- 192f0
		x"03304eb9", -- 192f4
		x"00004af4", -- 192f8
		x"08ac0000", -- 192fc
		x"00c14aac", -- 19300
		x"0048660e", -- 19304
		x"08380000", -- 19308
		x"fed26606", -- 1930c
		x"08ec0000", -- 19310
		x"00c141fa", -- 19314
		x"fca44a2c", -- 19318
		x"00a96604", -- 1931c
		x"41fafc80", -- 19320
		x"2f081f3c", -- 19324
		x"00011b7c", -- 19328
		x"0001ffef", -- 1932c
		x"486dffef", -- 19330
		x"4eba018a", -- 19334
		x"4e7548e7", -- 19338
		x"c0082878", -- 1933c
		x"fed408ec", -- 19340
		x"0005000a", -- 19344
		x"082c0006", -- 19348
		x"000a6618", -- 1934c
		x"4eb90000", -- 19350
		x"57e84eb9", -- 19354
		x"00005830", -- 19358
		x"7000322c", -- 1935c
		x"00565341", -- 19360
		x"4eac003c", -- 19364
		x"08ac0002", -- 19368
		x"000b6720", -- 1936c
		x"11ec00ca", -- 19370
		x"fdd2197c", -- 19374
		x"000300bb", -- 19378
		x"08ec0003", -- 1937c
		x"00c008ac", -- 19380
		x"000100c0", -- 19384
		x"670611ec", -- 19388
		x"00cbfdd2", -- 1938c
		x"297c0001", -- 19390
		x"8bc600c2", -- 19394
		x"297c0001", -- 19398
		x"8b1e00c6", -- 1939c
		x"197c0003", -- 193a0
		x"00ba08ec", -- 193a4
		x"000000c0", -- 193a8
		x"08ec0002", -- 193ac
		x"00c008ec", -- 193b0
		x"000700c0", -- 193b4
		x"4cdf1003", -- 193b8
		x"6000f808", -- 193bc
		x"2878fed4", -- 193c0
		x"297c2020", -- 193c4
		x"202000ca", -- 193c8
		x"297c0001", -- 193cc
		x"933a00c2", -- 193d0
		x"42ac00c6", -- 193d4
		x"422c00c1", -- 193d8
		x"47ec00ca", -- 193dc
		x"294b00b6", -- 193e0
		x"422c00ba", -- 193e4
		x"422c00bb", -- 193e8
		x"422c00c0", -- 193ec
		x"396c0046", -- 193f0
		x"00bc576c", -- 193f4
		x"00bc396c", -- 193f8
		x"005600be", -- 193fc
		x"08ec0007", -- 19400
		x"00c04e75", -- 19404
		x"205f2878", -- 19408
		x"fed44280", -- 1940c
		x"4281302c", -- 19410
		x"0046e240", -- 19414
		x"5240321f", -- 19418
		x"3b41fff4", -- 1941c
		x"4eac003c", -- 19420
		x"4ed0205f", -- 19424
		x"245f34ad", -- 19428
		x"fff44ed0", -- 1942c
		x"2878fed4", -- 19430
		x"302c0046", -- 19434
		x"e2405240", -- 19438
		x"3600322d", -- 1943c
		x"fff44eac", -- 19440
		x"003c1018", -- 19444
		x"67085243", -- 19448
		x"4eac0036", -- 1944c
		x"60f44e75", -- 19450
		x"2878fed4", -- 19454
		x"42804282", -- 19458
		x"302c0046", -- 1945c
		x"e2403400", -- 19460
		x"5240322d", -- 19464
		x"fff44eac", -- 19468
		x"003c5342", -- 1946c
		x"70204eac", -- 19470
		x"003651ca", -- 19474
		x"fff84e75", -- 19478
		x"2878fed4", -- 1947c
		x"42873e2c", -- 19480
		x"00565347", -- 19484
		x"60224286", -- 19488
		x"42804281", -- 1948c
		x"3c2c0046", -- 19490
		x"e2863006", -- 19494
		x"52403207", -- 19498
		x"4eac003c", -- 1949c
		x"53467020", -- 194a0
		x"4eac0036", -- 194a4
		x"51cefffa", -- 194a8
		x"be6dfff4", -- 194ac
		x"670451cf", -- 194b0
		x"ffd63f2d", -- 194b4
		x"fff44eba", -- 194b8
		x"ff4c4e75", -- 194bc
		x"205f225f", -- 194c0
		x"101f245f", -- 194c4
		x"2f084e56", -- 194c8
		x"ffe82d49", -- 194cc
		x"fff01d40", -- 194d0
		x"ffe82d4a", -- 194d4
		x"fffc422e", -- 194d8
		x"ffe9206e", -- 194dc
		x"fff04a10", -- 194e0
		x"670000ae", -- 194e4
		x"4a2effe8", -- 194e8
		x"670a3f3c", -- 194ec
		x"00014eba", -- 194f0
		x"ff146008", -- 194f4
		x"486effec", -- 194f8
		x"4ebaff28", -- 194fc
		x"6100ff7a", -- 19500
		x"42aefff4", -- 19504
		x"2d6efffc", -- 19508
		x"fff86700", -- 1950c
		x"0076206e", -- 19510
		x"fff8122c", -- 19514
		x"00c1c228", -- 19518
		x"0004b228", -- 1951c
		x"00046658", -- 19520
		x"10280005", -- 19524
		x"6d000052", -- 19528
		x"b07c0003", -- 1952c
		x"6e00004a", -- 19530
		x"e340323b", -- 19534
		x"00064efb", -- 19538
		x"1002003e", -- 1953c
		x"001a0008", -- 19540
		x"00382f2e", -- 19544
		x"fff8486e", -- 19548
		x"ffe92f2e", -- 1954c
		x"fff02268", -- 19550
		x"00064e91", -- 19554
		x"206efff8", -- 19558
		x"2d48fff4", -- 1955c
		x"41e8001a", -- 19560
		x"30106c04", -- 19564
		x"41f50000", -- 19568
		x"6100fec2", -- 1956c
		x"526dfff4", -- 19570
		x"600641e8", -- 19574
		x"000660e8", -- 19578
		x"206efff8", -- 1957c
		x"2d50fff8", -- 19580
		x"668c206e", -- 19584
		x"fff04210", -- 19588
		x"486effea", -- 1958c
		x"4ebafe94", -- 19590
		x"3f2effea", -- 19594
		x"4ebafe6e", -- 19598
		x"3600206e", -- 1959c
		x"fffc4a28", -- 195a0
		x"00056610", -- 195a4
		x"6100feaa", -- 195a8
		x"206efffc", -- 195ac
		x"41e80006", -- 195b0
		x"6100fe7a", -- 195b4
		x"2878fed4", -- 195b8
		x"396dfff4", -- 195bc
		x"00be3943", -- 195c0
		x"00bc197c", -- 195c4
		x"000300bb", -- 195c8
		x"08ec0003", -- 195cc
		x"00c008ec", -- 195d0
		x"000700c0", -- 195d4
		x"4eb90000", -- 195d8
		x"6d784a2c", -- 195dc
		x"00c06df4", -- 195e0
		x"526dfff4", -- 195e4
		x"202c00ca", -- 195e8
		x"103c0020", -- 195ec
		x"e0980c00", -- 195f0
		x"0020660a", -- 195f4
		x"e0980c00", -- 195f8
		x"00206602", -- 195fc
		x"e0982940", -- 19600
		x"00ca2d6e", -- 19604
		x"fffcfff8", -- 19608
		x"206efff8", -- 1960c
		x"122c00c1", -- 19610
		x"c2280004", -- 19614
		x"b2280004", -- 19618
		x"66161428", -- 1961c
		x"00050c02", -- 19620
		x"00026706", -- 19624
		x"0c020001", -- 19628
		x"6606b0a8", -- 1962c
		x"0016670e", -- 19630
		x"20502d48", -- 19634
		x"fff866d4", -- 19638
		x"2d6efff4", -- 1963c
		x"fff8206e", -- 19640
		x"fff82f08", -- 19644
		x"486effe9", -- 19648
		x"2f2efff0", -- 1964c
		x"20680006", -- 19650
		x"4e904a2e", -- 19654
		x"ffe96700", -- 19658
		x"fe824a2e", -- 1965c
		x"ffe8660c", -- 19660
		x"3f2effec", -- 19664
		x"6100fd9e", -- 19668
		x"6100fe0e", -- 1966c
		x"4e5e4e75", -- 19670
		x"205f141f", -- 19674
		x"121f245f", -- 19678
		x"225f7600", -- 1967c
		x"1612c602", -- 19680
		x"e22b1283", -- 19684
		x"4ed0205f", -- 19688
		x"141f121f", -- 1968c
		x"245f161f", -- 19690
		x"e32bc602", -- 19694
		x"18124602", -- 19698
		x"c8028803", -- 1969c
		x"14844ed0", -- 196a0
		x"205f101f", -- 196a4
		x"225f245f", -- 196a8
		x"42814282", -- 196ac
		x"42831211", -- 196b0
		x"54496016", -- 196b4
		x"16115449", -- 196b8
		x"1403e84a", -- 196bc
		x"0243000f", -- 196c0
		x"05006704", -- 196c4
		x"07d26002", -- 196c8
		x"079251c9", -- 196cc
		x"ffe84ed0", -- 196d0
		x"265f2e1f", -- 196d4
		x"285f2f0b", -- 196d8
		x"41f90040", -- 196dc
		x"800047f0", -- 196e0
		x"70007c00", -- 196e4
		x"1c1b6000", -- 196e8
		x"0076301b", -- 196ec
		x"0c00007e", -- 196f0
		x"66044614", -- 196f4
		x"60680c00", -- 196f8
		x"002b660c", -- 196fc
		x"321b0241", -- 19700
		x"00ffd314", -- 19704
		x"60000054", -- 19708
		x"0c00002a", -- 1970c
		x"6610030b", -- 19710
		x"0001584b", -- 19714
		x"14144882", -- 19718
		x"c5c11882", -- 1971c
		x"60380c00", -- 19720
		x"003c660e", -- 19724
		x"321b0241", -- 19728
		x"00ff1414", -- 1972c
		x"e32a1882", -- 19730
		x"60280c00", -- 19734
		x"003e660e", -- 19738
		x"321b0241", -- 1973c
		x"00ff1414", -- 19740
		x"e22a1882", -- 19744
		x"60140c00", -- 19748
		x"00416616", -- 1974c
		x"321b0241", -- 19750
		x"00ffc314", -- 19754
		x"60049c7c", -- 19758
		x"00019c7c", -- 1975c
		x"000151ce", -- 19760
		x"ff8a4e75", -- 19764
		x"4e75436f", -- 19768
		x"6e666967", -- 1976c
		x"75726520", -- 19770
		x"4d6f6465", -- 19774
		x"20466169", -- 19778
		x"6c656400", -- 1977c
		x"45455052", -- 19780
		x"4f4d2068", -- 19784
		x"61732062", -- 19788
		x"61642069", -- 1978c
		x"6e666f72", -- 19790
		x"6d617469", -- 19794
		x"6f6e0054", -- 19798
		x"6f6f206d", -- 1979c
		x"75636820", -- 197a0
		x"64617461", -- 197a4
		x"20746f20", -- 197a8
		x"73617665", -- 197ac
		x"00454550", -- 197b0
		x"524f4d20", -- 197b4
		x"4c6f6164", -- 197b8
		x"20736563", -- 197bc
		x"74696f6e", -- 197c0
		x"206d6973", -- 197c4
		x"73696e67", -- 197c8
		x"00454550", -- 197cc
		x"524f4d20", -- 197d0
		x"44656661", -- 197d4
		x"756c7473", -- 197d8
		x"20736563", -- 197dc
		x"74696f6e", -- 197e0
		x"206d6973", -- 197e4
		x"73696e67", -- 197e8
		x"00546f6f", -- 197ec
		x"206d616e", -- 197f0
		x"7920636f", -- 197f4
		x"6e666967", -- 197f8
		x"75726174", -- 197fc
		x"696f6e20", -- 19800
		x"73617665", -- 19804
		x"73004361", -- 19808
		x"6e206e6f", -- 1980c
		x"74207361", -- 19810
		x"76652063", -- 19814
		x"6f6e6669", -- 19818
		x"67757261", -- 1981c
		x"74696f6e", -- 19820
		x"00454550", -- 19824
		x"524f4d20", -- 19828
		x"63616e20", -- 1982c
		x"6e6f7420", -- 19830
		x"73617665", -- 19834
		x"20696e66", -- 19838
		x"6f726d61", -- 1983c
		x"74696f6e", -- 19840
		x"000048e7", -- 19844
		x"78807000", -- 19848
		x"72007603", -- 1984c
		x"78001218", -- 19850
		x"0c010020", -- 19854
		x"66064a44", -- 19858
		x"66246018", -- 1985c
		x"923c0030", -- 19860
		x"6d1c0c01", -- 19864
		x"00096e16", -- 19868
		x"d0802400", -- 1986c
		x"e580d082", -- 19870
		x"d0817801", -- 19874
		x"51cbffd8", -- 19878
		x"4cdf011e", -- 1987c
		x"4e7570ff", -- 19880
		x"60f648e7", -- 19884
		x"e08010fc", -- 19888
		x"002010fc", -- 1988c
		x"002010fc", -- 19890
		x"0020720a", -- 19894
		x"7430600c", -- 19898
		x"80c14840", -- 1989c
		x"d0421100", -- 198a0
		x"42404840", -- 198a4
		x"b08164f0", -- 198a8
		x"d0421100", -- 198ac
		x"4cdf0107", -- 198b0
		x"4e7513fc", -- 198b4
		x"00530040", -- 198b8
		x"000313fc", -- 198bc
		x"00cc0040", -- 198c0
		x"00050839", -- 198c4
		x"00040040", -- 198c8
		x"00034e75", -- 198cc
		x"08f80006", -- 198d0
		x"feda4dfa", -- 198d4
		x"001a4a39", -- 198d8
		x"00400001", -- 198dc
		x"66107208", -- 198e0
		x"b2390040", -- 198e4
		x"00056606", -- 198e8
		x"08b80006", -- 198ec
		x"feda4e75", -- 198f0
		x"4e56fff6", -- 198f4
		x"422efffb", -- 198f8
		x"2d7c0000", -- 198fc
		x"0001fffc", -- 19900
		x"206e000a", -- 19904
		x"202efffc", -- 19908
		x"10300800", -- 1990c
		x"b02e0008", -- 19910
		x"66081d7c", -- 19914
		x"0001fffb", -- 19918
		x"60580c00", -- 1991c
		x"00ff660c", -- 19920
		x"42aefffc", -- 19924
		x"1d7c0001", -- 19928
		x"fffb6046", -- 1992c
		x"202efffc", -- 19930
		x"5c802248", -- 19934
		x"222efffc", -- 19938
		x"58817400", -- 1993c
		x"14311800", -- 19940
		x"e1827200", -- 19944
		x"12300800", -- 19948
		x"d481e382", -- 1994c
		x"2d42fff6", -- 19950
		x"6f16d4ae", -- 19954
		x"fffc0c82", -- 19958
		x"00000fff", -- 1995c
		x"6c0a202e", -- 19960
		x"fff6d1ae", -- 19964
		x"fffc600a", -- 19968
		x"42aefffc", -- 1996c
		x"1d7c0001", -- 19970
		x"fffb4a2e", -- 19974
		x"fffb6788", -- 19978
		x"2d6efffc", -- 1997c
		x"000e4e5e", -- 19980
		x"205f5c4f", -- 19984
		x"4ed04e56", -- 19988
		x"fff6422e", -- 1998c
		x"ffff2d6e", -- 19990
		x"0008fff6", -- 19994
		x"06ae0000", -- 19998
		x"0014000c", -- 1999c
		x"206e0010", -- 199a0
		x"202e000c", -- 199a4
		x"4a300800", -- 199a8
		x"660c42ae", -- 199ac
		x"000c1d7c", -- 199b0
		x"0001ffff", -- 199b4
		x"604e202e", -- 199b8
		x"000c7201", -- 199bc
		x"b2300800", -- 199c0
		x"66425c80", -- 199c4
		x"10300800", -- 199c8
		x"b02efff6", -- 199cc
		x"6636202e", -- 199d0
		x"000c5080", -- 199d4
		x"10300800", -- 199d8
		x"b02efff7", -- 199dc
		x"6626700a", -- 199e0
		x"d0ae000c", -- 199e4
		x"10300800", -- 199e8
		x"b02efff8", -- 199ec
		x"6616700c", -- 199f0
		x"d0ae000c", -- 199f4
		x"10300800", -- 199f8
		x"b02efff9", -- 199fc
		x"66061d7c", -- 19a00
		x"0001ffff", -- 19a04
		x"4a2effff", -- 19a08
		x"6640206e", -- 19a0c
		x"0010202e", -- 19a10
		x"000c5480", -- 19a14
		x"72001230", -- 19a18
		x"0800e341", -- 19a1c
		x"48c12d41", -- 19a20
		x"fffa4aae", -- 19a24
		x"fffa6e08", -- 19a28
		x"3b7c0001", -- 19a2c
		x"fffe6032", -- 19a30
		x"202efffa", -- 19a34
		x"d1ae000c", -- 19a38
		x"0cae0000", -- 19a3c
		x"0fff000c", -- 19a40
		x"6f083b7c", -- 19a44
		x"0002fffe", -- 19a48
		x"60184a2e", -- 19a4c
		x"ffff6700", -- 19a50
		x"ff4c2d6e", -- 19a54
		x"000c0014", -- 19a58
		x"4e5e205f", -- 19a5c
		x"defc000c", -- 19a60
		x"4ed043fa", -- 19a64
		x"fd1841f8", -- 19a68
		x"fdd210d9", -- 19a6c
		x"66fc7000", -- 19a70
		x"302dfffe", -- 19a74
		x"53484eba", -- 19a78
		x"fe0a5648", -- 19a7c
		x"10bc0000", -- 19a80
		x"41f8fdd2", -- 19a84
		x"4efa23d0", -- 19a88
		x"4e56fffa", -- 19a8c
		x"102e0008", -- 19a90
		x"0200007f", -- 19a94
		x"1d400008", -- 19a98
		x"422effff", -- 19a9c
		x"06ae0000", -- 19aa0
		x"0014000a", -- 19aa4
		x"206e000e", -- 19aa8
		x"202e000a", -- 19aac
		x"4a300800", -- 19ab0
		x"660c42ae", -- 19ab4
		x"000a1d7c", -- 19ab8
		x"0001ffff", -- 19abc
		x"601e7201", -- 19ac0
		x"b2300800", -- 19ac4
		x"6616700e", -- 19ac8
		x"d0ae000a", -- 19acc
		x"10300800", -- 19ad0
		x"b02e0008", -- 19ad4
		x"66061d7c", -- 19ad8
		x"0001ffff", -- 19adc
		x"4a2effff", -- 19ae0
		x"6640206e", -- 19ae4
		x"000e202e", -- 19ae8
		x"000a5480", -- 19aec
		x"72001230", -- 19af0
		x"0800e341", -- 19af4
		x"48c12d41", -- 19af8
		x"fffa6e0a", -- 19afc
		x"3b7c0003", -- 19b00
		x"fffe6000", -- 19b04
		x"ff5e202e", -- 19b08
		x"fffad1ae", -- 19b0c
		x"000a0cae", -- 19b10
		x"00000fff", -- 19b14
		x"000a6f0a", -- 19b18
		x"3b7c0004", -- 19b1c
		x"fffe6000", -- 19b20
		x"ff424a2e", -- 19b24
		x"ffff6700", -- 19b28
		x"ff7c2d6e", -- 19b2c
		x"000a0012", -- 19b30
		x"4e5e205f", -- 19b34
		x"defc000a", -- 19b38
		x"4ed04e56", -- 19b3c
		x"fffc206e", -- 19b40
		x"000c226e", -- 19b44
		x"00082011", -- 19b48
		x"54807200", -- 19b4c
		x"12300800", -- 19b50
		x"e34148c1", -- 19b54
		x"2d41fffc", -- 19b58
		x"6e0a3b7c", -- 19b5c
		x"0005fffe", -- 19b60
		x"6000ff00", -- 19b64
		x"206e0008", -- 19b68
		x"202efffc", -- 19b6c
		x"d1904e5e", -- 19b70
		x"205f504f", -- 19b74
		x"4ed04e56", -- 19b78
		x"fff4206e", -- 19b7c
		x"00082d68", -- 19b80
		x"fff4fffc", -- 19b84
		x"22680008", -- 19b88
		x"2028fff0", -- 19b8c
		x"54807200", -- 19b90
		x"12310800", -- 19b94
		x"2141ffea", -- 19b98
		x"2028ffea", -- 19b9c
		x"91a8fff8", -- 19ba0
		x"6c0841fa", -- 19ba4
		x"fbf36000", -- 19ba8
		x"22ae7001", -- 19bac
		x"206e0008", -- 19bb0
		x"2d68ffea", -- 19bb4
		x"fff4b0ae", -- 19bb8
		x"fff46e2e", -- 19bbc
		x"2d40fff8", -- 19bc0
		x"206e0008", -- 19bc4
		x"22680008", -- 19bc8
		x"2028fff0", -- 19bcc
		x"2468000c", -- 19bd0
		x"2228fff4", -- 19bd4
		x"15b10800", -- 19bd8
		x"180054a8", -- 19bdc
		x"fff454a8", -- 19be0
		x"fff0202e", -- 19be4
		x"fff85280", -- 19be8
		x"68cc4aae", -- 19bec
		x"000c6700", -- 19bf0
		x"0084206e", -- 19bf4
		x"00082268", -- 19bf8
		x"000c202e", -- 19bfc
		x"fffc7201", -- 19c00
		x"b2310800", -- 19c04
		x"6600006e", -- 19c08
		x"7012d0ae", -- 19c0c
		x"fffc4a31", -- 19c10
		x"0800660c", -- 19c14
		x"7012d0ae", -- 19c18
		x"fffc13ae", -- 19c1c
		x"000f0800", -- 19c20
		x"206e0008", -- 19c24
		x"2268000c", -- 19c28
		x"202efffc", -- 19c2c
		x"50804a31", -- 19c30
		x"08006640", -- 19c34
		x"202efffc", -- 19c38
		x"5c804231", -- 19c3c
		x"0800202e", -- 19c40
		x"000c2268", -- 19c44
		x"000c222e", -- 19c48
		x"fffc5081", -- 19c4c
		x"45f90040", -- 19c50
		x"001013b2", -- 19c54
		x"08001800", -- 19c58
		x"2268000c", -- 19c5c
		x"700ad0ae", -- 19c60
		x"fffc4231", -- 19c64
		x"08002268", -- 19c68
		x"000c700c", -- 19c6c
		x"d0aefffc", -- 19c70
		x"42310800", -- 19c74
		x"206e0008", -- 19c78
		x"2028fff8", -- 19c7c
		x"6c06d0bc", -- 19c80
		x"000000ff", -- 19c84
		x"e0802268", -- 19c88
		x"000c720c", -- 19c8c
		x"d2adffde", -- 19c90
		x"13801800", -- 19c94
		x"2028fff8", -- 19c98
		x"02800000", -- 19c9c
		x"00ff2268", -- 19ca0
		x"000c720e", -- 19ca4
		x"d2adffde", -- 19ca8
		x"13801800", -- 19cac
		x"2268000c", -- 19cb0
		x"2028fff4", -- 19cb4
		x"42310800", -- 19cb8
		x"4e5e205f", -- 19cbc
		x"504f4ed0", -- 19cc0
		x"4e56ffdc", -- 19cc4
		x"70ff1200", -- 19cc8
		x"206e000c", -- 19ccc
		x"52801181", -- 19cd0
		x"08000c80", -- 19cd4
		x"00000fff", -- 19cd8
		x"6df2598f", -- 19cdc
		x"2f2e0008", -- 19ce0
		x"1f3c0001", -- 19ce4
		x"4ebafc0a", -- 19ce8
		x"2b5fffde", -- 19cec
		x"660841fa", -- 19cf0
		x"fabd6000", -- 19cf4
		x"2162206e", -- 19cf8
		x"0008202d", -- 19cfc
		x"ffde5c80", -- 19d00
		x"2248222d", -- 19d04
		x"ffde5881", -- 19d08
		x"74001431", -- 19d0c
		x"1800e182", -- 19d10
		x"72001230", -- 19d14
		x"0800d481", -- 19d18
		x"2d42fff8", -- 19d1c
		x"202efff8", -- 19d20
		x"e380d0ad", -- 19d24
		x"ffde5380", -- 19d28
		x"2b40ffe2", -- 19d2c
		x"206e0008", -- 19d30
		x"202dffde", -- 19d34
		x"226e000c", -- 19d38
		x"220013b0", -- 19d3c
		x"08001800", -- 19d40
		x"206e0008", -- 19d44
		x"202dffde", -- 19d48
		x"5480226e", -- 19d4c
		x"000c222d", -- 19d50
		x"ffde5481", -- 19d54
		x"13b00800", -- 19d58
		x"1800206e", -- 19d5c
		x"0008202d", -- 19d60
		x"ffde5880", -- 19d64
		x"226e000c", -- 19d68
		x"222dffde", -- 19d6c
		x"588113b0", -- 19d70
		x"08001800", -- 19d74
		x"206e0008", -- 19d78
		x"202dffde", -- 19d7c
		x"5c80226e", -- 19d80
		x"000c222d", -- 19d84
		x"ffde5c81", -- 19d88
		x"13b00800", -- 19d8c
		x"1800206e", -- 19d90
		x"0008202d", -- 19d94
		x"ffde5080", -- 19d98
		x"226e000c", -- 19d9c
		x"222dffde", -- 19da0
		x"508113b0", -- 19da4
		x"08001800", -- 19da8
		x"206e0008", -- 19dac
		x"700ad0ad", -- 19db0
		x"ffde226e", -- 19db4
		x"000c720a", -- 19db8
		x"d2adffde", -- 19dbc
		x"13b00800", -- 19dc0
		x"180004ae", -- 19dc4
		x"0000000a", -- 19dc8
		x"fff8202e", -- 19dcc
		x"fff86c06", -- 19dd0
		x"d0bc0000", -- 19dd4
		x"00ffe080", -- 19dd8
		x"206e000c", -- 19ddc
		x"720cd2ad", -- 19de0
		x"ffde1180", -- 19de4
		x"1800202e", -- 19de8
		x"fff80280", -- 19dec
		x"000000ff", -- 19df0
		x"206e000c", -- 19df4
		x"720ed2ad", -- 19df8
		x"ffde1180", -- 19dfc
		x"1800206e", -- 19e00
		x"00087010", -- 19e04
		x"d0adffde", -- 19e08
		x"226e000c", -- 19e0c
		x"7210d2ad", -- 19e10
		x"ffde13b0", -- 19e14
		x"08001800", -- 19e18
		x"206e0008", -- 19e1c
		x"7012d0ad", -- 19e20
		x"ffde226e", -- 19e24
		x"000c7212", -- 19e28
		x"d2adffde", -- 19e2c
		x"13b00800", -- 19e30
		x"18007014", -- 19e34
		x"d0adffde", -- 19e38
		x"2d40fff4", -- 19e3c
		x"206e000c", -- 19e40
		x"202efff4", -- 19e44
		x"42300800", -- 19e48
		x"2d6efff4", -- 19e4c
		x"fff0422e", -- 19e50
		x"ffef422e", -- 19e54
		x"ffe5206e", -- 19e58
		x"0008202e", -- 19e5c
		x"fff07200", -- 19e60
		x"12300800", -- 19e64
		x"6d0000c8", -- 19e68
		x"b27c0002", -- 19e6c
		x"6e0000c0", -- 19e70
		x"e341303b", -- 19e74
		x"10064efb", -- 19e78
		x"00020006", -- 19e7c
		x"001000ae", -- 19e80
		x"1d7c0001", -- 19e84
		x"ffef6000", -- 19e88
		x"00a6206e", -- 19e8c
		x"00087012", -- 19e90
		x"d0aefff0", -- 19e94
		x"72001230", -- 19e98
		x"08002d41", -- 19e9c
		x"ffe62f2d", -- 19ea0
		x"fff62f0e", -- 19ea4
		x"487a007a", -- 19ea8
		x"2b4ffff6", -- 19eac
		x"206e0008", -- 19eb0
		x"202efff0", -- 19eb4
		x"5080222e", -- 19eb8
		x"ffe643f9", -- 19ebc
		x"00400010", -- 19ec0
		x"12311800", -- 19ec4
		x"b2300800", -- 19ec8
		x"57c00200", -- 19ecc
		x"00011d40", -- 19ed0
		x"ffe56740", -- 19ed4
		x"202efff0", -- 19ed8
		x"d0bc0000", -- 19edc
		x"00104a30", -- 19ee0
		x"08006d30", -- 19ee4
		x"48415241", -- 19ee8
		x"22411011", -- 19eec
		x"08800007", -- 19ef0
		x"222efff0", -- 19ef4
		x"d2bc0000", -- 19ef8
		x"000eb030", -- 19efc
		x"10006714", -- 19f00
		x"222efff0", -- 19f04
		x"d2bc0000", -- 19f08
		x"0010b030", -- 19f0c
		x"10006704", -- 19f10
		x"42aeffe5", -- 19f14
		x"2b6f0008", -- 19f18
		x"fff6defc", -- 19f1c
		x"000c6006", -- 19f20
		x"2c5f2b5f", -- 19f24
		x"fff66006", -- 19f28
		x"1d7c0001", -- 19f2c
		x"ffe54a2e", -- 19f30
		x"ffef661c", -- 19f34
		x"4a2effe5", -- 19f38
		x"670a42a7", -- 19f3c
		x"2f0e4eba", -- 19f40
		x"fc36600c", -- 19f44
		x"2f2e0008", -- 19f48
		x"486efff0", -- 19f4c
		x"4ebafbec", -- 19f50
		x"0cae0000", -- 19f54
		x"0ffffff0", -- 19f58
		x"6f061d7c", -- 19f5c
		x"0001ffef", -- 19f60
		x"4a2effef", -- 19f64
		x"6700feec", -- 19f68
		x"598f2f2e", -- 19f6c
		x"00081f3c", -- 19f70
		x"00034eba", -- 19f74
		x"f97c2d5f", -- 19f78
		x"ffe06608", -- 19f7c
		x"41faf84b", -- 19f80
		x"60001ed4", -- 19f84
		x"422effef", -- 19f88
		x"2d7c0000", -- 19f8c
		x"0001ffe6", -- 19f90
		x"422effe5", -- 19f94
		x"42aeffdc", -- 19f98
		x"2f2dfff6", -- 19f9c
		x"2f0e487a", -- 19fa0
		x"008c2b4f", -- 19fa4
		x"fff6202e", -- 19fa8
		x"ffe641f9", -- 19fac
		x"00400010", -- 19fb0
		x"1d700800", -- 19fb4
		x"ffdd598f", -- 19fb8
		x"2f2e000c", -- 19fbc
		x"2f2dffde", -- 19fc0
		x"2f2effdc", -- 19fc4
		x"4ebaf9c0", -- 19fc8
		x"2d5ffff0", -- 19fcc
		x"6650598f", -- 19fd0
		x"2f2e0008", -- 19fd4
		x"2f2effe0", -- 19fd8
		x"2f2effdc", -- 19fdc
		x"4ebaf9a8", -- 19fe0
		x"2d5ffff0", -- 19fe4
		x"66327060", -- 19fe8
		x"b02effdd", -- 19fec
		x"62281d7c", -- 19ff0
		x"0001ffdf", -- 19ff4
		x"598f2f2e", -- 19ff8
		x"00082f2e", -- 19ffc
		x"ffe0206e", -- 1a000
		x"ffdc1f10", -- 1a004
		x"4ebafa82", -- 1a008
		x"2d5ffff0", -- 1a00c
		x"56c00200", -- 1a010
		x"00011d40", -- 1a014
		x"ffe56006", -- 1a018
		x"1d7c0001", -- 1a01c
		x"ffe52b6f", -- 1a020
		x"0008fff6", -- 1a024
		x"defc000c", -- 1a028
		x"4efa0008", -- 1a02c
		x"2c5f2b5f", -- 1a030
		x"fff64a2e", -- 1a034
		x"ffe5670a", -- 1a038
		x"2f2effe6", -- 1a03c
		x"2f0e4eba", -- 1a040
		x"fb3654ae", -- 1a044
		x"ffe67030", -- 1a048
		x"b0aeffe6", -- 1a04c
		x"6c061d7c", -- 1a050
		x"0001ffef", -- 1a054
		x"4a2effef", -- 1a058
		x"6700ff36", -- 1a05c
		x"2d6effe0", -- 1a060
		x"fff0422e", -- 1a064
		x"ffef422e", -- 1a068
		x"ffe5206e", -- 1a06c
		x"0008202e", -- 1a070
		x"fff07200", -- 1a074
		x"12300800", -- 1a078
		x"6d72b27c", -- 1a07c
		x"00026e6c", -- 1a080
		x"e341303b", -- 1a084
		x"10064efb", -- 1a088
		x"00020006", -- 1a08c
		x"000c000e", -- 1a090
		x"1d7c0001", -- 1a094
		x"ffef6054", -- 1a098
		x"206e000c", -- 1a09c
		x"202efff0", -- 1a0a0
		x"5c801d70", -- 1a0a4
		x"0800ffdc", -- 1a0a8
		x"202efff0", -- 1a0ac
		x"50801d70", -- 1a0b0
		x"0800ffdd", -- 1a0b4
		x"700ad0ae", -- 1a0b8
		x"fff01d70", -- 1a0bc
		x"0800ffde", -- 1a0c0
		x"700cd0ae", -- 1a0c4
		x"fff01d70", -- 1a0c8
		x"0800ffdf", -- 1a0cc
		x"598f2f2e", -- 1a0d0
		x"000c2f2d", -- 1a0d4
		x"ffde2f2e", -- 1a0d8
		x"ffdc4eba", -- 1a0dc
		x"f8aa2d5f", -- 1a0e0
		x"fffc57c0", -- 1a0e4
		x"02000001", -- 1a0e8
		x"1d40ffe5", -- 1a0ec
		x"4a2effe5", -- 1a0f0
		x"670a42a7", -- 1a0f4
		x"2f0e4eba", -- 1a0f8
		x"fa7e600c", -- 1a0fc
		x"2f2e0008", -- 1a100
		x"486efff0", -- 1a104
		x"4ebafa34", -- 1a108
		x"0cae0000", -- 1a10c
		x"0ffffff0", -- 1a110
		x"6f061d7c", -- 1a114
		x"0001ffef", -- 1a118
		x"4a2effef", -- 1a11c
		x"6700ff48", -- 1a120
		x"4e5e205f", -- 1a124
		x"504f4ed0", -- 1a128
		x"4e56fffa", -- 1a12c
		x"42ae0012", -- 1a130
		x"422effff", -- 1a134
		x"06ae0000", -- 1a138
		x"0014000a", -- 1a13c
		x"206e000e", -- 1a140
		x"202e000a", -- 1a144
		x"10300800", -- 1a148
		x"b02e0008", -- 1a14c
		x"660e1d7c", -- 1a150
		x"0001ffff", -- 1a154
		x"2d6e000a", -- 1a158
		x"0012604a", -- 1a15c
		x"202e000a", -- 1a160
		x"4a300800", -- 1a164
		x"66081d7c", -- 1a168
		x"0001ffff", -- 1a16c
		x"6038202e", -- 1a170
		x"000a5480", -- 1a174
		x"72001230", -- 1a178
		x"0800e341", -- 1a17c
		x"48c12d41", -- 1a180
		x"fffa6608", -- 1a184
		x"1d7c0001", -- 1a188
		x"ffff601a", -- 1a18c
		x"202efffa", -- 1a190
		x"d1ae000a", -- 1a194
		x"0cae0000", -- 1a198
		x"0fff000a", -- 1a19c
		x"5ec00200", -- 1a1a0
		x"00011d40", -- 1a1a4
		x"ffff4a2e", -- 1a1a8
		x"ffff6790", -- 1a1ac
		x"4e5e205f", -- 1a1b0
		x"defc000a", -- 1a1b4
		x"4ed02f2f", -- 1a1b8
		x"00082f3c", -- 1a1bc
		x"00000030", -- 1a1c0
		x"4eb90000", -- 1a1c4
		x"0ae4245f", -- 1a1c8
		x"225f205f", -- 1a1cc
		x"205042a8", -- 1a1d0
		x"00004228", -- 1a1d4
		x"0004117c", -- 1a1d8
		x"00030005", -- 1a1dc
		x"41e80006", -- 1a1e0
		x"10d966fc", -- 1a1e4
		x"4ed22f2f", -- 1a1e8
		x"000c2f3c", -- 1a1ec
		x"00000036", -- 1a1f0
		x"4eb90000", -- 1a1f4
		x"0ae4285f", -- 1a1f8
		x"2e1f265f", -- 1a1fc
		x"205f2050", -- 1a200
		x"42a80000", -- 1a204
		x"42280004", -- 1a208
		x"117c0001", -- 1a20c
		x"0005117c", -- 1a210
		x"00200016", -- 1a214
		x"11530017", -- 1a218
		x"116b0001", -- 1a21c
		x"0018116b", -- 1a220
		x"00020019", -- 1a224
		x"45e8001a", -- 1a228
		x"14db66fc", -- 1a22c
		x"21470006", -- 1a230
		x"42a8000a", -- 1a234
		x"42a8000e", -- 1a238
		x"42a80012", -- 1a23c
		x"4ed441f9", -- 1a240
		x"00018e16", -- 1a244
		x"2e884e56", -- 1a248
		x"ffd82d6d", -- 1a24c
		x"ffdefff4", -- 1a250
		x"42aefff8", -- 1a254
		x"202efff4", -- 1a258
		x"b0adffe2", -- 1a25c
		x"6e2c4aae", -- 1a260
		x"fff86626", -- 1a264
		x"41f90040", -- 1a268
		x"8000226d", -- 1a26c
		x"fff02200", -- 1a270
		x"12311800", -- 1a274
		x"b2300800", -- 1a278
		x"660654ae", -- 1a27c
		x"fff46008", -- 1a280
		x"2d7c0000", -- 1a284
		x"0001fff8", -- 1a288
		x"60ca4aae", -- 1a28c
		x"fff86f00", -- 1a290
		x"02082d6d", -- 1a294
		x"ffdefff4", -- 1a298
		x"206dfff0", -- 1a29c
		x"7012d0ae", -- 1a2a0
		x"fff42248", -- 1a2a4
		x"7210d2ae", -- 1a2a8
		x"fff47400", -- 1a2ac
		x"14311800", -- 1a2b0
		x"e1827200", -- 1a2b4
		x"12300800", -- 1a2b8
		x"d4812d42", -- 1a2bc
		x"fff80cae", -- 1a2c0
		x"0000ffff", -- 1a2c4
		x"fff8660c", -- 1a2c8
		x"41faf51f", -- 1a2cc
		x"4eb90000", -- 1a2d0
		x"57cc6038", -- 1a2d4
		x"52aefff8", -- 1a2d8
		x"202efff8", -- 1a2dc
		x"6c06d0bc", -- 1a2e0
		x"000000ff", -- 1a2e4
		x"e080206d", -- 1a2e8
		x"fff07210", -- 1a2ec
		x"d2aefff4", -- 1a2f0
		x"11801800", -- 1a2f4
		x"202efff8", -- 1a2f8
		x"02800000", -- 1a2fc
		x"00ff206d", -- 1a300
		x"fff07212", -- 1a304
		x"d2aefff4", -- 1a308
		x"11801800", -- 1a30c
		x"206dfff0", -- 1a310
		x"202efff4", -- 1a314
		x"5c802248", -- 1a318
		x"222efff4", -- 1a31c
		x"58817400", -- 1a320
		x"14311800", -- 1a324
		x"e1827200", -- 1a328
		x"12300800", -- 1a32c
		x"d4812d42", -- 1a330
		x"fffc6f00", -- 1a334
		x"0098202e", -- 1a338
		x"fffc0280", -- 1a33c
		x"00000003", -- 1a340
		x"6600008a", -- 1a344
		x"082e0000", -- 1a348
		x"ffff670e", -- 1a34c
		x"3b7c0000", -- 1a350
		x"fffe41fa", -- 1a354
		x"f4b26000", -- 1a358
		x"1afe206d", -- 1a35c
		x"fff0700a", -- 1a360
		x"d0aefff4", -- 1a364
		x"2248222e", -- 1a368
		x"fff45081", -- 1a36c
		x"74001431", -- 1a370
		x"1800e182", -- 1a374
		x"72001230", -- 1a378
		x"0800d481", -- 1a37c
		x"2d42ffe2", -- 1a380
		x"206dfff0", -- 1a384
		x"202efff4", -- 1a388
		x"50804230", -- 1a38c
		x"0800206d", -- 1a390
		x"fff0700a", -- 1a394
		x"d0aefff4", -- 1a398
		x"42300800", -- 1a39c
		x"206dfff0", -- 1a3a0
		x"202efff4", -- 1a3a4
		x"538041f0", -- 1a3a8
		x"0800282e", -- 1a3ac
		x"fffce384", -- 1a3b0
		x"4eb90000", -- 1a3b4
		x"4eaa5343", -- 1a3b8
		x"4643206d", -- 1a3bc
		x"fff0202e", -- 1a3c0
		x"fff45080", -- 1a3c4
		x"43f00800", -- 1a3c8
		x"07890000", -- 1a3cc
		x"3b7c0001", -- 1a3d0
		x"fffe4eba", -- 1a3d4
		x"f4de6700", -- 1a3d8
		x"ff7a42ae", -- 1a3dc
		x"fff82d6d", -- 1a3e0
		x"ffdefff4", -- 1a3e4
		x"202efff4", -- 1a3e8
		x"b0adffe2", -- 1a3ec
		x"6e00008e", -- 1a3f0
		x"206dfff0", -- 1a3f4
		x"1d700800", -- 1a3f8
		x"ffeb202e", -- 1a3fc
		x"fff441f9", -- 1a400
		x"00408000", -- 1a404
		x"122effeb", -- 1a408
		x"b2300800", -- 1a40c
		x"6766202e", -- 1a410
		x"fff441f9", -- 1a414
		x"00408000", -- 1a418
		x"11aeffeb", -- 1a41c
		x"08004eb9", -- 1a420
		x"000051d8", -- 1a424
		x"2d40ffec", -- 1a428
		x"90bc0000", -- 1a42c
		x"09c42d40", -- 1a430
		x"fff0202e", -- 1a434
		x"fff441f9", -- 1a438
		x"00408000", -- 1a43c
		x"122effeb", -- 1a440
		x"b2300800", -- 1a444
		x"670e4eb9", -- 1a448
		x"000051d8", -- 1a44c
		x"b0aefff0", -- 1a450
		x"6d0260de", -- 1a454
		x"202efff4", -- 1a458
		x"41f90040", -- 1a45c
		x"8000122e", -- 1a460
		x"ffebb230", -- 1a464
		x"08006708", -- 1a468
		x"41faf3b7", -- 1a46c
		x"600019e8", -- 1a470
		x"52aefff8", -- 1a474
		x"54aefff4", -- 1a478
		x"6000ff6a", -- 1a47c
		x"13fc0000", -- 1a480
		x"00400001", -- 1a484
		x"08390004", -- 1a488
		x"00400003", -- 1a48c
		x"670a3b7c", -- 1a490
		x"0002fffe", -- 1a494
		x"6000febc", -- 1a498
		x"4e5e205f", -- 1a49c
		x"defc000c", -- 1a4a0
		x"4ed04e56", -- 1a4a4
		x"fff4202d", -- 1a4a8
		x"ffde5c80", -- 1a4ac
		x"41f90040", -- 1a4b0
		x"8000222d", -- 1a4b4
		x"ffde5881", -- 1a4b8
		x"43f90040", -- 1a4bc
		x"80007400", -- 1a4c0
		x"14311800", -- 1a4c4
		x"e1827200", -- 1a4c8
		x"12300800", -- 1a4cc
		x"d4812d42", -- 1a4d0
		x"fff804ae", -- 1a4d4
		x"0000000a", -- 1a4d8
		x"fff8202e", -- 1a4dc
		x"fff86c06", -- 1a4e0
		x"d0bc0000", -- 1a4e4
		x"00ffe080", -- 1a4e8
		x"206dfff0", -- 1a4ec
		x"720cd2ad", -- 1a4f0
		x"ffde1180", -- 1a4f4
		x"1800202e", -- 1a4f8
		x"fff80280", -- 1a4fc
		x"000000ff", -- 1a500
		x"720ed2ad", -- 1a504
		x"ffde1180", -- 1a508
		x"18007014", -- 1a50c
		x"d0adffde", -- 1a510
		x"42300800", -- 1a514
		x"7015d0ad", -- 1a518
		x"ffde2d6d", -- 1a51c
		x"ffe2fff4", -- 1a520
		x"b0aefff4", -- 1a524
		x"6e1a2d40", -- 1a528
		x"fffc206d", -- 1a52c
		x"fff0202e", -- 1a530
		x"fffc11bc", -- 1a534
		x"00ff0800", -- 1a538
		x"202efffc", -- 1a53c
		x"528068e0", -- 1a540
		x"2f2e0010", -- 1a544
		x"2f2e000c", -- 1a548
		x"2f2e0008", -- 1a54c
		x"4ebafcf8", -- 1a550
		x"41fa000e", -- 1a554
		x"4eb90000", -- 1a558
		x"57cc4ef9", -- 1a55c
		x"00004bf4", -- 1a560
		x"4d757374", -- 1a564
		x"20637963", -- 1a568
		x"6c652053", -- 1a56c
		x"50552070", -- 1a570
		x"6f776572", -- 1a574
		x"20746f20", -- 1a578
		x"636f6d70", -- 1a57c
		x"6c657465", -- 1a580
		x"20646566", -- 1a584
		x"61756c74", -- 1a588
		x"20736574", -- 1a58c
		x"75700000", -- 1a590
		x"4e560000", -- 1a594
		x"4e5e205f", -- 1a598
		x"defc000c", -- 1a59c
		x"4ed04e56", -- 1a5a0
		x"0000206e", -- 1a5a4
		x"000c10bc", -- 1a5a8
		x"00014e5e", -- 1a5ac
		x"205fdefc", -- 1a5b0
		x"000c4ed0", -- 1a5b4
		x"285f205f", -- 1a5b8
		x"221f2e8c", -- 1a5bc
		x"50817000", -- 1a5c0
		x"226dfff0", -- 1a5c4
		x"10311800", -- 1a5c8
		x"907c0060", -- 1a5cc
		x"48c04eba", -- 1a5d0
		x"f2b2117c", -- 1a5d4
		x"00000003", -- 1a5d8
		x"4e752078", -- 1a5dc
		x"fed42068", -- 1a5e0
		x"00b60c28", -- 1a5e4
		x"00200003", -- 1a5e8
		x"4e754e56", -- 1a5ec
		x"fff4206e", -- 1a5f0
		x"000c4210", -- 1a5f4
		x"206e0008", -- 1a5f8
		x"42104eba", -- 1a5fc
		x"ffde660c", -- 1a600
		x"206e000c", -- 1a604
		x"10bc0001", -- 1a608
		x"600000a0", -- 1a60c
		x"2078fed4", -- 1a610
		x"206800b6", -- 1a614
		x"4ebaf22c", -- 1a618
		x"2d40fffc", -- 1a61c
		x"206e0010", -- 1a620
		x"20280012", -- 1a624
		x"5c8041f9", -- 1a628
		x"00408000", -- 1a62c
		x"122effff", -- 1a630
		x"b2300800", -- 1a634
		x"6574206e", -- 1a638
		x"00102028", -- 1a63c
		x"00125080", -- 1a640
		x"41f90040", -- 1a644
		x"8000b230", -- 1a648
		x"0800625e", -- 1a64c
		x"206dfff0", -- 1a650
		x"226e0010", -- 1a654
		x"2029000e", -- 1a658
		x"50807200", -- 1a65c
		x"12300800", -- 1a660
		x"70609240", -- 1a664
		x"48c12d41", -- 1a668
		x"fff8202e", -- 1a66c
		x"fffc242d", -- 1a670
		x"ffdab081", -- 1a674
		x"672c0102", -- 1a678
		x"66300382", -- 1a67c
		x"01c22b42", -- 1a680
		x"ffda7060", -- 1a684
		x"d0aefffc", -- 1a688
		x"206dfff0", -- 1a68c
		x"226e0010", -- 1a690
		x"2229000e", -- 1a694
		x"50811180", -- 1a698
		x"1800206e", -- 1a69c
		x"000810bc", -- 1a6a0
		x"0001206e", -- 1a6a4
		x"000c10bc", -- 1a6a8
		x"00014e5e", -- 1a6ac
		x"205fdefc", -- 1a6b0
		x"000c4ed0", -- 1a6b4
		x"4e56ffd4", -- 1a6b8
		x"206e000c", -- 1a6bc
		x"4210206e", -- 1a6c0
		x"00084a10", -- 1a6c4
		x"6728206e", -- 1a6c8
		x"00102f28", -- 1a6cc
		x"00122f28", -- 1a6d0
		x"000e486e", -- 1a6d4
		x"fffc4eba", -- 1a6d8
		x"fedc41ee", -- 1a6dc
		x"fffc226e", -- 1a6e0
		x"001043e9", -- 1a6e4
		x"003112d8", -- 1a6e8
		x"66fc6000", -- 1a6ec
		x"01f8206d", -- 1a6f0
		x"fff0226e", -- 1a6f4
		x"00102029", -- 1a6f8
		x"000e5080", -- 1a6fc
		x"72001230", -- 1a700
		x"08007060", -- 1a704
		x"924048c1", -- 1a708
		x"2d41ffe8", -- 1a70c
		x"206e0010", -- 1a710
		x"20280012", -- 1a714
		x"5c807200", -- 1a718
		x"43f90040", -- 1a71c
		x"80001231", -- 1a720
		x"08002d41", -- 1a724
		x"ffec1231", -- 1a728
		x"08022d41", -- 1a72c
		x"fff02d68", -- 1a730
		x"000affdc", -- 1a734
		x"66000068", -- 1a738
		x"486effdc", -- 1a73c
		x"2f3c0000", -- 1a740
		x"00304eb9", -- 1a744
		x"00000ae4", -- 1a748
		x"2d6effdc", -- 1a74c
		x"ffd8206e", -- 1a750
		x"ffd842a8", -- 1a754
		x"00004228", -- 1a758
		x"0004117c", -- 1a75c
		x"00000005", -- 1a760
		x"43e80006", -- 1a764
		x"45fa018a", -- 1a768
		x"12da66fc", -- 1a76c
		x"4eba01ca", -- 1a770
		x"284841ec", -- 1a774
		x"000a202e", -- 1a778
		x"ffec4eba", -- 1a77c
		x"f10641ec", -- 1a780
		x"000f202e", -- 1a784
		x"fff04eba", -- 1a788
		x"f0fa486e", -- 1a78c
		x"ffe0487a", -- 1a790
		x"015e4eba", -- 1a794
		x"fa22206e", -- 1a798
		x"ffdc20ae", -- 1a79c
		x"ffe0206e", -- 1a7a0
		x"00104aa8", -- 1a7a4
		x"000a663e", -- 1a7a8
		x"486effe4", -- 1a7ac
		x"4868001a", -- 1a7b0
		x"487afe38", -- 1a7b4
		x"4ebafa30", -- 1a7b8
		x"2d6effe4", -- 1a7bc
		x"ffd8206e", -- 1a7c0
		x"ffd842a8", -- 1a7c4
		x"000a226e", -- 1a7c8
		x"00102169", -- 1a7cc
		x"000e000e", -- 1a7d0
		x"21690012", -- 1a7d4
		x"0012206e", -- 1a7d8
		x"ffe020ae", -- 1a7dc
		x"ffe42d6e", -- 1a7e0
		x"ffe4ffe0", -- 1a7e4
		x"6022206e", -- 1a7e8
		x"ffdc2068", -- 1a7ec
		x"00002d68", -- 1a7f0
		x"0000ffe4", -- 1a7f4
		x"206e0010", -- 1a7f8
		x"43e8001a", -- 1a7fc
		x"246effe4", -- 1a800
		x"41ea001a", -- 1a804
		x"10d966fc", -- 1a808
		x"206e0010", -- 1a80c
		x"4aa8000a", -- 1a810
		x"6644486e", -- 1a814
		x"ffe4487a", -- 1a818
		x"00f14eba", -- 1a81c
		x"f99a206e", -- 1a820
		x"ffe020ae", -- 1a824
		x"ffe42d6e", -- 1a828
		x"ffe4ffe0", -- 1a82c
		x"486effe4", -- 1a830
		x"2f3c0000", -- 1a834
		x"00304eb9", -- 1a838
		x"00000ae4", -- 1a83c
		x"2d6effe4", -- 1a840
		x"ffd8206e", -- 1a844
		x"ffd842a8", -- 1a848
		x"00004228", -- 1a84c
		x"0004117c", -- 1a850
		x"00030005", -- 1a854
		x"600e206e", -- 1a858
		x"ffe42068", -- 1a85c
		x"00002d68", -- 1a860
		x"0000ffe4", -- 1a864
		x"2d6effe4", -- 1a868
		x"ffd8202e", -- 1a86c
		x"ffec2d6e", -- 1a870
		x"fff0ffd4", -- 1a874
		x"286effd8", -- 1a878
		x"49ec0006", -- 1a87c
		x"b0aeffd4", -- 1a880
		x"6e262d40", -- 1a884
		x"fff4b0ae", -- 1a888
		x"ffe86714", -- 1a88c
		x"222dffda", -- 1a890
		x"0101670c", -- 1a894
		x"204c4eba", -- 1a898
		x"efea564c", -- 1a89c
		x"18bc0000", -- 1a8a0
		x"202efff4", -- 1a8a4
		x"528068d4", -- 1a8a8
		x"206e0010", -- 1a8ac
		x"4aa8000a", -- 1a8b0
		x"661a206e", -- 1a8b4
		x"ffe0216e", -- 1a8b8
		x"ffe40000", -- 1a8bc
		x"2d6effe4", -- 1a8c0
		x"ffe0206e", -- 1a8c4
		x"0010216e", -- 1a8c8
		x"ffdc000a", -- 1a8cc
		x"206e0008", -- 1a8d0
		x"10bc0001", -- 1a8d4
		x"2f2effdc", -- 1a8d8
		x"42272f2e", -- 1a8dc
		x"00084eb9", -- 1a8e0
		x"000194c0", -- 1a8e4
		x"4e5e205f", -- 1a8e8
		x"defc000c", -- 1a8ec
		x"4ed02000", -- 1a8f0
		x"54797065", -- 1a8f4
		x"2020202e", -- 1a8f8
		x"2e202020", -- 1a8fc
		x"20657863", -- 1a900
		x"65707420", -- 1a904
		x"75736564", -- 1a908
		x"00202075", -- 1a90c
		x"73656420", -- 1a910
		x"73656c65", -- 1a914
		x"63742063", -- 1a918
		x"6f646573", -- 1a91c
		x"20617265", -- 1a920
		x"3a002052", -- 1a924
		x"45545552", -- 1a928
		x"4e203f20", -- 1a92c
		x"0020454e", -- 1a930
		x"54455220", -- 1a934
		x"3f200000", -- 1a938
		x"48e70088", -- 1a93c
		x"534941fa", -- 1a940
		x"ffe22878", -- 1a944
		x"fed44a2c", -- 1a948
		x"00a96604", -- 1a94c
		x"41faffdf", -- 1a950
		x"12d866fc", -- 1a954
		x"4cdf1100", -- 1a958
		x"4e754e56", -- 1a95c
		x"fff642ae", -- 1a960
		x"0010422e", -- 1a964
		x"ffff422e", -- 1a968
		x"fffe42ae", -- 1a96c
		x"fffa206d", -- 1a970
		x"fff0202e", -- 1a974
		x"000c5880", -- 1a978
		x"72001230", -- 1a97c
		x"0800e341", -- 1a980
		x"48c1d2ae", -- 1a984
		x"000c5581", -- 1a988
		x"2d41000c", -- 1a98c
		x"54ae000c", -- 1a990
		x"206dfff0", -- 1a994
		x"202e000c", -- 1a998
		x"72001230", -- 1a99c
		x"08006d00", -- 1a9a0
		x"00fcb27c", -- 1a9a4
		x"00096e00", -- 1a9a8
		x"00f4e341", -- 1a9ac
		x"303b1006", -- 1a9b0
		x"4efb0002", -- 1a9b4
		x"0014001e", -- 1a9b8
		x"00380066", -- 1a9bc
		x"007e00d0", -- 1a9c0
		x"00e600e6", -- 1a9c4
		x"00660066", -- 1a9c8
		x"1d7c0001", -- 1a9cc
		x"ffff6000", -- 1a9d0
		x"00d654ae", -- 1a9d4
		x"000c206d", -- 1a9d8
		x"fff0202e", -- 1a9dc
		x"000c7200", -- 1a9e0
		x"12300800", -- 1a9e4
		x"2d41fffa", -- 1a9e8
		x"600000bc", -- 1a9ec
		x"206dfff0", -- 1a9f0
		x"202e000c", -- 1a9f4
		x"58802248", -- 1a9f8
		x"222e000c", -- 1a9fc
		x"54817400", -- 1aa00
		x"14311800", -- 1aa04
		x"e1827200", -- 1aa08
		x"12300800", -- 1aa0c
		x"d4812d42", -- 1aa10
		x"fffa58ae", -- 1aa14
		x"000c6000", -- 1aa18
		x"008e54ae", -- 1aa1c
		x"000c202e", -- 1aa20
		x"fffab0ae", -- 1aa24
		x"000857c0", -- 1aa28
		x"02000001", -- 1aa2c
		x"1d40fffe", -- 1aa30
		x"607454ae", -- 1aa34
		x"000c206d", -- 1aa38
		x"fff0202e", -- 1aa3c
		x"000c7200", -- 1aa40
		x"12300800", -- 1aa44
		x"2d41fff6", -- 1aa48
		x"202efffa", -- 1aa4c
		x"b0ae0008", -- 1aa50
		x"6d26202e", -- 1aa54
		x"0008d0ae", -- 1aa58
		x"fff6b0ae", -- 1aa5c
		x"fffa6f18", -- 1aa60
		x"202efffa", -- 1aa64
		x"90ae0008", -- 1aa68
		x"5280e380", -- 1aa6c
		x"d1ae000c", -- 1aa70
		x"1d7c0001", -- 1aa74
		x"fffe600a", -- 1aa78
		x"202efff6", -- 1aa7c
		x"e380d1ae", -- 1aa80
		x"000c6022", -- 1aa84
		x"58ae000c", -- 1aa88
		x"202efffa", -- 1aa8c
		x"b0ae0008", -- 1aa90
		x"57c00200", -- 1aa94
		x"00011d40", -- 1aa98
		x"fffe600a", -- 1aa9c
		x"3b7c0006", -- 1aaa0
		x"fffe6000", -- 1aaa4
		x"efbe102e", -- 1aaa8
		x"ffff660a", -- 1aaac
		x"102efffe", -- 1aab0
		x"66046000", -- 1aab4
		x"fed84a2e", -- 1aab8
		x"fffe6706", -- 1aabc
		x"2d6e000c", -- 1aac0
		x"00104e5e", -- 1aac4
		x"205f504f", -- 1aac8
		x"4ed04e56", -- 1aacc
		x"fffa41fa", -- 1aad0
		x"00b2246e", -- 1aad4
		x"000843d2", -- 1aad8
		x"12d866fc", -- 1aadc
		x"700cd0ae", -- 1aae0
		x"001041f9", -- 1aae4
		x"00408000", -- 1aae8
		x"720ad2ae", -- 1aaec
		x"001043f9", -- 1aaf0
		x"00408000", -- 1aaf4
		x"74001431", -- 1aaf8
		x"1800e182", -- 1aafc
		x"72001230", -- 1ab00
		x"0800d481", -- 1ab04
		x"2d42fffc", -- 1ab08
		x"598f2f2e", -- 1ab0c
		x"000c2f2e", -- 1ab10
		x"fffc4eba", -- 1ab14
		x"fe462d5f", -- 1ab18
		x"fffc6f5c", -- 1ab1c
		x"486efffb", -- 1ab20
		x"206dfff0", -- 1ab24
		x"202efffc", -- 1ab28
		x"48700800", -- 1ab2c
		x"700ed0ae", -- 1ab30
		x"001041f9", -- 1ab34
		x"00408000", -- 1ab38
		x"1f300800", -- 1ab3c
		x"7010d0ae", -- 1ab40
		x"001041f9", -- 1ab44
		x"00408000", -- 1ab48
		x"1f300800", -- 1ab4c
		x"4eb90001", -- 1ab50
		x"9674486e", -- 1ab54
		x"fffb7012", -- 1ab58
		x"d0ae0010", -- 1ab5c
		x"2f004eb9", -- 1ab60
		x"000196d4", -- 1ab64
		x"7000102e", -- 1ab68
		x"fffb206e", -- 1ab6c
		x"00084eba", -- 1ab70
		x"ed12117c", -- 1ab74
		x"00000003", -- 1ab78
		x"4e5e205f", -- 1ab7c
		x"defc000c", -- 1ab80
		x"4ed06e6e", -- 1ab84
		x"6e004e56", -- 1ab88
		x"ffee206e", -- 1ab8c
		x"000c4210", -- 1ab90
		x"206e0008", -- 1ab94
		x"42104eba", -- 1ab98
		x"fa42660c", -- 1ab9c
		x"206e000c", -- 1aba0
		x"10bc0001", -- 1aba4
		x"60000160", -- 1aba8
		x"2078fed4", -- 1abac
		x"206800b6", -- 1abb0
		x"4ebaec90", -- 1abb4
		x"2d40fff4", -- 1abb8
		x"6d00014c", -- 1abbc
		x"0c800000", -- 1abc0
		x"00ff6e00", -- 1abc4
		x"01421d6e", -- 1abc8
		x"fff7ffef", -- 1abcc
		x"206e0010", -- 1abd0
		x"2d680012", -- 1abd4
		x"fff8700c", -- 1abd8
		x"d0aefff8", -- 1abdc
		x"41f90040", -- 1abe0
		x"8000720a", -- 1abe4
		x"d2aefff8", -- 1abe8
		x"43f90040", -- 1abec
		x"80007400", -- 1abf0
		x"14311800", -- 1abf4
		x"e1827200", -- 1abf8
		x"12300800", -- 1abfc
		x"d4812d42", -- 1ac00
		x"fff4598f", -- 1ac04
		x"206e0010", -- 1ac08
		x"2f28000e", -- 1ac0c
		x"2f2efff4", -- 1ac10
		x"4ebafd48", -- 1ac14
		x"2d5ffff4", -- 1ac18
		x"660a3b7c", -- 1ac1c
		x"0007fffe", -- 1ac20
		x"6000ee40", -- 1ac24
		x"202efff8", -- 1ac28
		x"5c8041f9", -- 1ac2c
		x"00408000", -- 1ac30
		x"122effef", -- 1ac34
		x"b2300800", -- 1ac38
		x"650000cc", -- 1ac3c
		x"202efff8", -- 1ac40
		x"508041f9", -- 1ac44
		x"00408000", -- 1ac48
		x"b2300800", -- 1ac4c
		x"620000b8", -- 1ac50
		x"7012d0ae", -- 1ac54
		x"fff841f9", -- 1ac58
		x"00408000", -- 1ac5c
		x"72001230", -- 1ac60
		x"0800e341", -- 1ac64
		x"48c1d2ae", -- 1ac68
		x"fff87014", -- 1ac6c
		x"d2802d41", -- 1ac70
		x"fffc486e", -- 1ac74
		x"ffef2f2e", -- 1ac78
		x"fffc4eb9", -- 1ac7c
		x"000196d4", -- 1ac80
		x"1f2effef", -- 1ac84
		x"206dfff0", -- 1ac88
		x"202efff4", -- 1ac8c
		x"48700800", -- 1ac90
		x"700ed0ae", -- 1ac94
		x"fff841f9", -- 1ac98
		x"00408000", -- 1ac9c
		x"1f300800", -- 1aca0
		x"7010d0ae", -- 1aca4
		x"fff841f9", -- 1aca8
		x"00408000", -- 1acac
		x"1f300800", -- 1acb0
		x"4eb90001", -- 1acb4
		x"968a206d", -- 1acb8
		x"fff0226e", -- 1acbc
		x"0010700e", -- 1acc0
		x"d0a90018", -- 1acc4
		x"48700800", -- 1acc8
		x"202efffc", -- 1accc
		x"41f90040", -- 1acd0
		x"80007200", -- 1acd4
		x"12300800", -- 1acd8
		x"e34148c1", -- 1acdc
		x"d2aefffc", -- 1ace0
		x"548141f9", -- 1ace4
		x"00408000", -- 1ace8
		x"48701800", -- 1acec
		x"1f2effef", -- 1acf0
		x"4eb90001", -- 1acf4
		x"96a4206e", -- 1acf8
		x"000c10bc", -- 1acfc
		x"0001206e", -- 1ad00
		x"000810bc", -- 1ad04
		x"00014e5e", -- 1ad08
		x"205fdefc", -- 1ad0c
		x"000c4ed0", -- 1ad10
		x"4e56ffe0", -- 1ad14
		x"206e000c", -- 1ad18
		x"4210206e", -- 1ad1c
		x"00084a10", -- 1ad20
		x"6728206e", -- 1ad24
		x"00102f28", -- 1ad28
		x"00122f28", -- 1ad2c
		x"000e486e", -- 1ad30
		x"fffc4eba", -- 1ad34
		x"fd9641ee", -- 1ad38
		x"fffc226e", -- 1ad3c
		x"001043e9", -- 1ad40
		x"003112d8", -- 1ad44
		x"66fc6000", -- 1ad48
		x"012a206e", -- 1ad4c
		x"00102d68", -- 1ad50
		x"000affe4", -- 1ad54
		x"660000e2", -- 1ad58
		x"486effe4", -- 1ad5c
		x"2f3c0000", -- 1ad60
		x"00304eb9", -- 1ad64
		x"00000ae4", -- 1ad68
		x"206effe4", -- 1ad6c
		x"2d48ffe0", -- 1ad70
		x"42a80000", -- 1ad74
		x"42280004", -- 1ad78
		x"117c0000", -- 1ad7c
		x"0005226e", -- 1ad80
		x"00102029", -- 1ad84
		x"00125c80", -- 1ad88
		x"720043f9", -- 1ad8c
		x"00408000", -- 1ad90
		x"12310800", -- 1ad94
		x"2d41fff0", -- 1ad98
		x"226e0010", -- 1ad9c
		x"20290012", -- 1ada0
		x"50807200", -- 1ada4
		x"43f90040", -- 1ada8
		x"80001231", -- 1adac
		x"08002d41", -- 1adb0
		x"fff443fa", -- 1adb4
		x"00ca45e8", -- 1adb8
		x"000614d9", -- 1adbc
		x"66fc224a", -- 1adc0
		x"4ebafb76", -- 1adc4
		x"284841ec", -- 1adc8
		x"000a202e", -- 1adcc
		x"fff04eba", -- 1add0
		x"eab241ec", -- 1add4
		x"000f202e", -- 1add8
		x"fff44eba", -- 1addc
		x"eaa6486e", -- 1ade0
		x"ffe8487a", -- 1ade4
		x"00984eba", -- 1ade8
		x"f3ce206e", -- 1adec
		x"ffe4216e", -- 1adf0
		x"ffe80000", -- 1adf4
		x"486effec", -- 1adf8
		x"206e0010", -- 1adfc
		x"4868001a", -- 1ae00
		x"487afd84", -- 1ae04
		x"4ebaf3e0", -- 1ae08
		x"2d6effec", -- 1ae0c
		x"ffe0206e", -- 1ae10
		x"ffe042a8", -- 1ae14
		x"000a226e", -- 1ae18
		x"00102169", -- 1ae1c
		x"000e000e", -- 1ae20
		x"21690012", -- 1ae24
		x"0012206e", -- 1ae28
		x"ffe8216e", -- 1ae2c
		x"ffec0000", -- 1ae30
		x"2d6effec", -- 1ae34
		x"ffe86022", -- 1ae38
		x"206effe4", -- 1ae3c
		x"20680000", -- 1ae40
		x"2d680000", -- 1ae44
		x"ffec206e", -- 1ae48
		x"001043e8", -- 1ae4c
		x"001a246e", -- 1ae50
		x"ffec41ea", -- 1ae54
		x"001a10d9", -- 1ae58
		x"66fc206e", -- 1ae5c
		x"000810bc", -- 1ae60
		x"00012f2e", -- 1ae64
		x"ffe44227", -- 1ae68
		x"2f2e0008", -- 1ae6c
		x"4eb90001", -- 1ae70
		x"94c04e5e", -- 1ae74
		x"205fdefc", -- 1ae78
		x"000c4ed0", -- 1ae7c
		x"20005479", -- 1ae80
		x"70652020", -- 1ae84
		x"202e2e20", -- 1ae88
		x"20200000", -- 1ae8c
		x"4e560000", -- 1ae90
		x"42ae0012", -- 1ae94
		x"58ae000a", -- 1ae98
		x"206e000e", -- 1ae9c
		x"202e000a", -- 1aea0
		x"4a300800", -- 1aea4
		x"67361030", -- 1aea8
		x"0800b02e", -- 1aeac
		x"00086608", -- 1aeb0
		x"2d6e000a", -- 1aeb4
		x"00126024", -- 1aeb8
		x"206e000e", -- 1aebc
		x"202e000a", -- 1aec0
		x"54807200", -- 1aec4
		x"12300800", -- 1aec8
		x"e54148c1", -- 1aecc
		x"e381202e", -- 1aed0
		x"000a5880", -- 1aed4
		x"d0812d40", -- 1aed8
		x"000a60bc", -- 1aedc
		x"4e5e205f", -- 1aee0
		x"defc000a", -- 1aee4
		x"4ed04e56", -- 1aee8
		x"fffc42ae", -- 1aeec
		x"0012206e", -- 1aef0
		x"000e202e", -- 1aef4
		x"000a5480", -- 1aef8
		x"72001230", -- 1aefc
		x"08002d41", -- 1af00
		x"fffc58ae", -- 1af04
		x"000a4aae", -- 1af08
		x"fffc6f24", -- 1af0c
		x"206e000e", -- 1af10
		x"202e000a", -- 1af14
		x"10300800", -- 1af18
		x"b02e0008", -- 1af1c
		x"66082d6e", -- 1af20
		x"000a0012", -- 1af24
		x"600a53ae", -- 1af28
		x"fffc50ae", -- 1af2c
		x"000a60d6", -- 1af30
		x"4e5e205f", -- 1af34
		x"defc000a", -- 1af38
		x"4ed04e56", -- 1af3c
		x"fffc42ae", -- 1af40
		x"0014206e", -- 1af44
		x"0010202e", -- 1af48
		x"000c5480", -- 1af4c
		x"72001230", -- 1af50
		x"08002d41", -- 1af54
		x"fffc58ae", -- 1af58
		x"000c4aae", -- 1af5c
		x"fffc6f46", -- 1af60
		x"206e0010", -- 1af64
		x"202e000c", -- 1af68
		x"54801030", -- 1af6c
		x"0800b02e", -- 1af70
		x"00096628", -- 1af74
		x"202e000c", -- 1af78
		x"58801030", -- 1af7c
		x"0800b02e", -- 1af80
		x"000a6618", -- 1af84
		x"202e000c", -- 1af88
		x"5c801030", -- 1af8c
		x"0800b02e", -- 1af90
		x"000b6608", -- 1af94
		x"2d6e000c", -- 1af98
		x"0014600a", -- 1af9c
		x"53aefffc", -- 1afa0
		x"50ae000c", -- 1afa4
		x"60b44e5e", -- 1afa8
		x"205fdefc", -- 1afac
		x"000c4ed0", -- 1afb0
		x"4e56fffa", -- 1afb4
		x"41fa011e", -- 1afb8
		x"246e0008", -- 1afbc
		x"43d212d8", -- 1afc0
		x"66fc202e", -- 1afc4
		x"00105080", -- 1afc8
		x"41f90040", -- 1afcc
		x"8000222e", -- 1afd0
		x"00105c81", -- 1afd4
		x"43f90040", -- 1afd8
		x"80007400", -- 1afdc
		x"14311800", -- 1afe0
		x"e1827200", -- 1afe4
		x"12300800", -- 1afe8
		x"d4812d42", -- 1afec
		x"fffc598f", -- 1aff0
		x"2f2e000c", -- 1aff4
		x"2f2efffc", -- 1aff8
		x"4ebaf960", -- 1affc
		x"2d5ffffc", -- 1b000
		x"6f0000c8", -- 1b004
		x"486efffb", -- 1b008
		x"206dfff0", -- 1b00c
		x"202efffc", -- 1b010
		x"48700800", -- 1b014
		x"700ad0ae", -- 1b018
		x"001041f9", -- 1b01c
		x"00408000", -- 1b020
		x"1f300800", -- 1b024
		x"700cd0ae", -- 1b028
		x"001041f9", -- 1b02c
		x"00408000", -- 1b030
		x"1f300800", -- 1b034
		x"4eb90001", -- 1b038
		x"9674598f", -- 1b03c
		x"48790040", -- 1b040
		x"80001f3c", -- 1b044
		x"00024eba", -- 1b048
		x"e8a82d5f", -- 1b04c
		x"fffc6f7a", -- 1b050
		x"598f4879", -- 1b054
		x"00408000", -- 1b058
		x"2f2efffc", -- 1b05c
		x"1f3c0003", -- 1b060
		x"4ebaf0c6", -- 1b064
		x"2d5ffffc", -- 1b068
		x"6f60598f", -- 1b06c
		x"48790040", -- 1b070
		x"80002f2e", -- 1b074
		x"fffc700e", -- 1b078
		x"d0ae0010", -- 1b07c
		x"41f90040", -- 1b080
		x"80001f30", -- 1b084
		x"08004eba", -- 1b088
		x"fe042d5f", -- 1b08c
		x"fffc6f3a", -- 1b090
		x"598f4879", -- 1b094
		x"00408000", -- 1b098
		x"2f2efffc", -- 1b09c
		x"1f2efffb", -- 1b0a0
		x"4ebafe44", -- 1b0a4
		x"2d5ffffc", -- 1b0a8
		x"6f20202e", -- 1b0ac
		x"fffc43f9", -- 1b0b0
		x"00408000", -- 1b0b4
		x"43f10800", -- 1b0b8
		x"206e0008", -- 1b0bc
		x"10e90002", -- 1b0c0
		x"10e90004", -- 1b0c4
		x"10e90006", -- 1b0c8
		x"42104e5e", -- 1b0cc
		x"205fdefc", -- 1b0d0
		x"000c4ed0", -- 1b0d4
		x"61616100", -- 1b0d8
		x"4e56fff4", -- 1b0dc
		x"206e000c", -- 1b0e0
		x"42104eba", -- 1b0e4
		x"f4f6660c", -- 1b0e8
		x"206e000c", -- 1b0ec
		x"10bc0001", -- 1b0f0
		x"60000156", -- 1b0f4
		x"206e0010", -- 1b0f8
		x"2d680012", -- 1b0fc
		x"fff4202e", -- 1b100
		x"fff45080", -- 1b104
		x"41f90040", -- 1b108
		x"8000222e", -- 1b10c
		x"fff45c81", -- 1b110
		x"43f90040", -- 1b114
		x"80007400", -- 1b118
		x"14311800", -- 1b11c
		x"e1827200", -- 1b120
		x"12300800", -- 1b124
		x"d4812d42", -- 1b128
		x"fffc598f", -- 1b12c
		x"206e0010", -- 1b130
		x"2f28000e", -- 1b134
		x"2f2efffc", -- 1b138
		x"4ebaf820", -- 1b13c
		x"2d5ffff8", -- 1b140
		x"6f000106", -- 1b144
		x"598f4879", -- 1b148
		x"00408000", -- 1b14c
		x"1f3c0002", -- 1b150
		x"4ebae79e", -- 1b154
		x"2d5ffffc", -- 1b158
		x"6f0000ee", -- 1b15c
		x"598f4879", -- 1b160
		x"00408000", -- 1b164
		x"2f2efffc", -- 1b168
		x"1f3c0003", -- 1b16c
		x"4ebaefba", -- 1b170
		x"2d5ffffc", -- 1b174
		x"6f0000d2", -- 1b178
		x"598f4879", -- 1b17c
		x"00408000", -- 1b180
		x"2f2efffc", -- 1b184
		x"700ed0ae", -- 1b188
		x"fff441f9", -- 1b18c
		x"00408000", -- 1b190
		x"1f300800", -- 1b194
		x"4ebafcf6", -- 1b198
		x"2d5ffffc", -- 1b19c
		x"6f0000aa", -- 1b1a0
		x"598f4879", -- 1b1a4
		x"00408000", -- 1b1a8
		x"2f2efffc", -- 1b1ac
		x"2078fed4", -- 1b1b0
		x"206800b6", -- 1b1b4
		x"2f104eba", -- 1b1b8
		x"fd822d5f", -- 1b1bc
		x"fffc6f00", -- 1b1c0
		x"0088202e", -- 1b1c4
		x"fffc41f9", -- 1b1c8
		x"00408000", -- 1b1cc
		x"1f300800", -- 1b1d0
		x"206dfff0", -- 1b1d4
		x"202efff8", -- 1b1d8
		x"48700800", -- 1b1dc
		x"700ad0ae", -- 1b1e0
		x"fff441f9", -- 1b1e4
		x"00408000", -- 1b1e8
		x"1f300800", -- 1b1ec
		x"700cd0ae", -- 1b1f0
		x"fff441f9", -- 1b1f4
		x"00408000", -- 1b1f8
		x"1f300800", -- 1b1fc
		x"4eb90001", -- 1b200
		x"968a206d", -- 1b204
		x"fff0226e", -- 1b208
		x"0010700e", -- 1b20c
		x"d0a9000e", -- 1b210
		x"48700800", -- 1b214
		x"7010d0ae", -- 1b218
		x"fff441f9", -- 1b21c
		x"00408000", -- 1b220
		x"48700800", -- 1b224
		x"202efffc", -- 1b228
		x"41f90040", -- 1b22c
		x"80001f30", -- 1b230
		x"08004eb9", -- 1b234
		x"000196a4", -- 1b238
		x"206e000c", -- 1b23c
		x"10bc0001", -- 1b240
		x"206e0008", -- 1b244
		x"10bc0001", -- 1b248
		x"4e5e205f", -- 1b24c
		x"defc000c", -- 1b250
		x"4ed04e56", -- 1b254
		x"fedc206e", -- 1b258
		x"000c4210", -- 1b25c
		x"206e0008", -- 1b260
		x"4a106728", -- 1b264
		x"206e0010", -- 1b268
		x"2f280012", -- 1b26c
		x"2f28000e", -- 1b270
		x"486efffc", -- 1b274
		x"4ebafd3a", -- 1b278
		x"41eefffc", -- 1b27c
		x"226e0010", -- 1b280
		x"43e90031", -- 1b284
		x"12d866fc", -- 1b288
		x"600001dc", -- 1b28c
		x"206e0010", -- 1b290
		x"2d68000a", -- 1b294
		x"fff46600", -- 1b298
		x"0194486e", -- 1b29c
		x"fff42f3c", -- 1b2a0
		x"00000030", -- 1b2a4
		x"4eb90000", -- 1b2a8
		x"0ae42d6e", -- 1b2ac
		x"fff4ffe0", -- 1b2b0
		x"206effe0", -- 1b2b4
		x"42a80000", -- 1b2b8
		x"42280004", -- 1b2bc
		x"117c0000", -- 1b2c0
		x"000543fa", -- 1b2c4
		x"01ae45e8", -- 1b2c8
		x"000614d9", -- 1b2cc
		x"66fc538a", -- 1b2d0
		x"2d4afedc", -- 1b2d4
		x"598f4879", -- 1b2d8
		x"00408000", -- 1b2dc
		x"1f3c0002", -- 1b2e0
		x"4ebae60e", -- 1b2e4
		x"2d5fffe8", -- 1b2e8
		x"6f0000d8", -- 1b2ec
		x"598f4879", -- 1b2f0
		x"00408000", -- 1b2f4
		x"2f2effe8", -- 1b2f8
		x"1f3c0003", -- 1b2fc
		x"4ebaee2a", -- 1b300
		x"2d5fffe8", -- 1b304
		x"6f0000bc", -- 1b308
		x"598f4879", -- 1b30c
		x"00408000", -- 1b310
		x"2f2effe8", -- 1b314
		x"206e0010", -- 1b318
		x"700ed0a8", -- 1b31c
		x"001241f9", -- 1b320
		x"00408000", -- 1b324
		x"1f300800", -- 1b328
		x"4ebafb62", -- 1b32c
		x"2d5fffe8", -- 1b330
		x"6f000090", -- 1b334
		x"202effe8", -- 1b338
		x"54807200", -- 1b33c
		x"41f90040", -- 1b340
		x"80001230", -- 1b344
		x"08002d41", -- 1b348
		x"ffec58ae", -- 1b34c
		x"ffe854ae", -- 1b350
		x"ffe8202e", -- 1b354
		x"ffe849f0", -- 1b358
		x"0800226e", -- 1b35c
		x"fedc7202", -- 1b360
		x"10140c00", -- 1b364
		x"00206702", -- 1b368
		x"12c0548c", -- 1b36c
		x"51c9fff2", -- 1b370
		x"42115cae", -- 1b374
		x"ffe82d49", -- 1b378
		x"fedc7002", -- 1b37c
		x"b0aeffec", -- 1b380
		x"6c16226e", -- 1b384
		x"fedc12fc", -- 1b388
		x"002c12fc", -- 1b38c
		x"002012bc", -- 1b390
		x"00002d49", -- 1b394
		x"fedc6024", -- 1b398
		x"7002b0ae", -- 1b39c
		x"ffec661c", -- 1b3a0
		x"226efedc", -- 1b3a4
		x"12fc0020", -- 1b3a8
		x"12fc006f", -- 1b3ac
		x"12fc0072", -- 1b3b0
		x"12fc0020", -- 1b3b4
		x"12bc0000", -- 1b3b8
		x"2d49fedc", -- 1b3bc
		x"53aeffec", -- 1b3c0
		x"668c226e", -- 1b3c4
		x"fedc5249", -- 1b3c8
		x"6100f56e", -- 1b3cc
		x"486efff8", -- 1b3d0
		x"487a009e", -- 1b3d4
		x"4ebaede0", -- 1b3d8
		x"206efff4", -- 1b3dc
		x"20aefff8", -- 1b3e0
		x"486efff0", -- 1b3e4
		x"206e0010", -- 1b3e8
		x"4868001a", -- 1b3ec
		x"487afcea", -- 1b3f0
		x"4ebaedf4", -- 1b3f4
		x"2d6efff0", -- 1b3f8
		x"ffe0206e", -- 1b3fc
		x"ffe042a8", -- 1b400
		x"000a226e", -- 1b404
		x"00102169", -- 1b408
		x"000e000e", -- 1b40c
		x"21690012", -- 1b410
		x"0012206e", -- 1b414
		x"fff820ae", -- 1b418
		x"fff02d6e", -- 1b41c
		x"fff0fff8", -- 1b420
		x"206e0010", -- 1b424
		x"216efff4", -- 1b428
		x"000a6022", -- 1b42c
		x"206efff4", -- 1b430
		x"20680000", -- 1b434
		x"2d680000", -- 1b438
		x"fff0206e", -- 1b43c
		x"001043e8", -- 1b440
		x"001a246e", -- 1b444
		x"fff041ea", -- 1b448
		x"001a10d9", -- 1b44c
		x"66fc206e", -- 1b450
		x"000810bc", -- 1b454
		x"00012f2e", -- 1b458
		x"fff44227", -- 1b45c
		x"2f2e0008", -- 1b460
		x"4eb90001", -- 1b464
		x"94c04e5e", -- 1b468
		x"205fdefc", -- 1b46c
		x"000c4ed0", -- 1b470
		x"20005479", -- 1b474
		x"70652000", -- 1b478
		x"4e56fffe", -- 1b47c
		x"42ae0012", -- 1b480
		x"422effff", -- 1b484
		x"58ae000a", -- 1b488
		x"206e000e", -- 1b48c
		x"202e000a", -- 1b490
		x"10300800", -- 1b494
		x"b02e0008", -- 1b498
		x"660e1d7c", -- 1b49c
		x"0001ffff", -- 1b4a0
		x"2d6e000a", -- 1b4a4
		x"00126028", -- 1b4a8
		x"206e000e", -- 1b4ac
		x"202e000a", -- 1b4b0
		x"4a300800", -- 1b4b4
		x"66081d7c", -- 1b4b8
		x"0001ffff", -- 1b4bc
		x"601254ae", -- 1b4c0
		x"000a206e", -- 1b4c4
		x"000e202e", -- 1b4c8
		x"000a4a30", -- 1b4cc
		x"080066ee", -- 1b4d0
		x"54ae000a", -- 1b4d4
		x"4a2effff", -- 1b4d8
		x"67ae4e5e", -- 1b4dc
		x"205fdefc", -- 1b4e0
		x"000a4ed0", -- 1b4e4
		x"285f265f", -- 1b4e8
		x"201f245f", -- 1b4ec
		x"45f20802", -- 1b4f0
		x"16d26704", -- 1b4f4
		x"548a60f8", -- 1b4f8
		x"4ed44e56", -- 1b4fc
		x"fff2246e", -- 1b500
		x"000843d2", -- 1b504
		x"4211202e", -- 1b508
		x"001041f9", -- 1b50c
		x"00408000", -- 1b510
		x"1d700800", -- 1b514
		x"fff32d7c", -- 1b518
		x"00408000", -- 1b51c
		x"fff4598f", -- 1b520
		x"2f2efff4", -- 1b524
		x"1f3c0002", -- 1b528
		x"4ebae3c6", -- 1b52c
		x"2d5ffff8", -- 1b530
		x"6f40598f", -- 1b534
		x"2f2efff4", -- 1b538
		x"2f2efff8", -- 1b53c
		x"1f3c0002", -- 1b540
		x"4ebaebe6", -- 1b544
		x"2d5ffffc", -- 1b548
		x"6f28598f", -- 1b54c
		x"2f2efff4", -- 1b550
		x"2f2efffc", -- 1b554
		x"1f2efff3", -- 1b558
		x"4ebaff1e", -- 1b55c
		x"2d5ffffc", -- 1b560
		x"6f102f2e", -- 1b564
		x"fff42f2e", -- 1b568
		x"fffc2f2e", -- 1b56c
		x"00084eba", -- 1b570
		x"ff744e5e", -- 1b574
		x"205fdefc", -- 1b578
		x"000c4ed0", -- 1b57c
		x"4e56fecc", -- 1b580
		x"206e0008", -- 1b584
		x"4a106734", -- 1b588
		x"2d6e0010", -- 1b58c
		x"ffc8206d", -- 1b590
		x"fff0226e", -- 1b594
		x"ffc82029", -- 1b598
		x"000e5080", -- 1b59c
		x"72001230", -- 1b5a0
		x"08007060", -- 1b5a4
		x"924048c1", -- 1b5a8
		x"2d41fffc", -- 1b5ac
		x"41e90031", -- 1b5b0
		x"202efffc", -- 1b5b4
		x"4ebae2cc", -- 1b5b8
		x"600002b2", -- 1b5bc
		x"206e0010", -- 1b5c0
		x"2d68000a", -- 1b5c4
		x"ffec6600", -- 1b5c8
		x"0282486e", -- 1b5cc
		x"ffec2f3c", -- 1b5d0
		x"00000030", -- 1b5d4
		x"4eb90000", -- 1b5d8
		x"0ae42d6e", -- 1b5dc
		x"ffecffc8", -- 1b5e0
		x"206effc8", -- 1b5e4
		x"42a80000", -- 1b5e8
		x"42280004", -- 1b5ec
		x"117c0000", -- 1b5f0
		x"000543fa", -- 1b5f4
		x"080045e8", -- 1b5f8
		x"000614d9", -- 1b5fc
		x"66fc224a", -- 1b600
		x"4ebaf336", -- 1b604
		x"41eefecc", -- 1b608
		x"700410fc", -- 1b60c
		x"002051c8", -- 1b610
		x"fffa226e", -- 1b614
		x"001043e9", -- 1b618
		x"001f700f", -- 1b61c
		x"10d951c8", -- 1b620
		x"fffc4210", -- 1b624
		x"486efff0", -- 1b628
		x"486efecc", -- 1b62c
		x"4ebaeb88", -- 1b630
		x"206effec", -- 1b634
		x"20aefff0", -- 1b638
		x"486effe8", -- 1b63c
		x"487a0249", -- 1b640
		x"4ebaeb74", -- 1b644
		x"206efff0", -- 1b648
		x"20aeffe8", -- 1b64c
		x"2d6effe8", -- 1b650
		x"fff0486e", -- 1b654
		x"ffe8487a", -- 1b658
		x"07184eba", -- 1b65c
		x"eb5a206e", -- 1b660
		x"fff020ae", -- 1b664
		x"ffe82d6e", -- 1b668
		x"ffe8fff0", -- 1b66c
		x"42aefff4", -- 1b670
		x"206e0010", -- 1b674
		x"20280012", -- 1b678
		x"5c802d40", -- 1b67c
		x"fffc202e", -- 1b680
		x"fffc41f9", -- 1b684
		x"00408000", -- 1b688
		x"4a300800", -- 1b68c
		x"660a1d7c", -- 1b690
		x"0001ffd1", -- 1b694
		x"6000014c", -- 1b698
		x"52aefff4", -- 1b69c
		x"486effe8", -- 1b6a0
		x"2f3c0000", -- 1b6a4
		x"00364eb9", -- 1b6a8
		x"00000ae4", -- 1b6ac
		x"246effe8", -- 1b6b0
		x"2d4affc8", -- 1b6b4
		x"43ea001a", -- 1b6b8
		x"701a12fc", -- 1b6bc
		x"002051c8", -- 1b6c0
		x"fffa12bc", -- 1b6c4
		x"00002f2e", -- 1b6c8
		x"fffc206e", -- 1b6cc
		x"00102f28", -- 1b6d0
		x"000e486e", -- 1b6d4
		x"ffd64eba", -- 1b6d8
		x"fe22202e", -- 1b6dc
		x"fff4206e", -- 1b6e0
		x"ffc841e8", -- 1b6e4
		x"001a4eba", -- 1b6e8
		x"e19a5688", -- 1b6ec
		x"10fc0020", -- 1b6f0
		x"10fc0020", -- 1b6f4
		x"43eeffd6", -- 1b6f8
		x"10d966fc", -- 1b6fc
		x"534810bc", -- 1b700
		x"0020206e", -- 1b704
		x"ffc842a8", -- 1b708
		x"00004228", -- 1b70c
		x"0004117c", -- 1b710
		x"00020005", -- 1b714
		x"42a8000a", -- 1b718
		x"226e0010", -- 1b71c
		x"2169000e", -- 1b720
		x"000e216e", -- 1b724
		x"fffc0012", -- 1b728
		x"117c0020", -- 1b72c
		x"00161168", -- 1b730
		x"001a0017", -- 1b734
		x"1168001b", -- 1b738
		x"00181168", -- 1b73c
		x"001c0019", -- 1b740
		x"202efffc", -- 1b744
		x"588043f9", -- 1b748
		x"00408000", -- 1b74c
		x"72001231", -- 1b750
		x"08005341", -- 1b754
		x"6d34b27c", -- 1b758
		x"00026e2e", -- 1b75c
		x"e341303b", -- 1b760
		x"10064efb", -- 1b764
		x"00020006", -- 1b768
		x"0010001a", -- 1b76c
		x"217c0001", -- 1b770
		x"a6b80006", -- 1b774
		x"601e217c", -- 1b778
		x"0001ad14", -- 1b77c
		x"00066014", -- 1b780
		x"217c0001", -- 1b784
		x"b2560006", -- 1b788
		x"600a3b7c", -- 1b78c
		x"0008fffe", -- 1b790
		x"6000e2d0", -- 1b794
		x"206efff0", -- 1b798
		x"216effe8", -- 1b79c
		x"00002d6e", -- 1b7a0
		x"ffe8fff0", -- 1b7a4
		x"202efffc", -- 1b7a8
		x"548041f9", -- 1b7ac
		x"00408000", -- 1b7b0
		x"72001230", -- 1b7b4
		x"0800e341", -- 1b7b8
		x"48c12d41", -- 1b7bc
		x"ffcc6e08", -- 1b7c0
		x"1d7c0001", -- 1b7c4
		x"ffd1601a", -- 1b7c8
		x"202effcc", -- 1b7cc
		x"d1aefffc", -- 1b7d0
		x"0cae0000", -- 1b7d4
		x"0ffffffc", -- 1b7d8
		x"5ec00200", -- 1b7dc
		x"00011d40", -- 1b7e0
		x"ffd14a2e", -- 1b7e4
		x"ffd16700", -- 1b7e8
		x"fe96486e", -- 1b7ec
		x"ffe8487a", -- 1b7f0
		x"00864eba", -- 1b7f4
		x"e9c2206e", -- 1b7f8
		x"fff020ae", -- 1b7fc
		x"ffe82d6e", -- 1b800
		x"ffe8fff0", -- 1b804
		x"486effe8", -- 1b808
		x"487a006e", -- 1b80c
		x"487aed90", -- 1b810
		x"4ebae9d4", -- 1b814
		x"206efff0", -- 1b818
		x"20aeffe8", -- 1b81c
		x"2d6effe8", -- 1b820
		x"fff0486e", -- 1b824
		x"ffe8487a", -- 1b828
		x"0548487a", -- 1b82c
		x"ed644eba", -- 1b830
		x"e9b6206e", -- 1b834
		x"fff020ae", -- 1b838
		x"ffe82d6e", -- 1b83c
		x"ffe8fff0", -- 1b840
		x"206e0010", -- 1b844
		x"216effec", -- 1b848
		x"000a206e", -- 1b84c
		x"000810bc", -- 1b850
		x"00012f2e", -- 1b854
		x"ffec1f3c", -- 1b858
		x"00012f2e", -- 1b85c
		x"00084eb9", -- 1b860
		x"000194c0", -- 1b864
		x"206e0008", -- 1b868
		x"10bc0001", -- 1b86c
		x"4e5e205f", -- 1b870
		x"defc000c", -- 1b874
		x"4ed02000", -- 1b878
		x"20205820", -- 1b87c
		x"20655869", -- 1b880
		x"74206d65", -- 1b884
		x"6e75006b", -- 1b888
		x"65797320", -- 1b88c
		x"46656174", -- 1b890
		x"75726520", -- 1b894
		x"20202020", -- 1b898
		x"20202020", -- 1b89c
		x"56616c75", -- 1b8a0
		x"65004e56", -- 1b8a4
		x"fffa42ae", -- 1b8a8
		x"0012422e", -- 1b8ac
		x"ffff58ae", -- 1b8b0
		x"000a206e", -- 1b8b4
		x"000e202e", -- 1b8b8
		x"000a1030", -- 1b8bc
		x"0800b02e", -- 1b8c0
		x"0008660e", -- 1b8c4
		x"2d6e000a", -- 1b8c8
		x"00121d7c", -- 1b8cc
		x"0001ffff", -- 1b8d0
		x"6052206e", -- 1b8d4
		x"000e202e", -- 1b8d8
		x"000a4a30", -- 1b8dc
		x"08006608", -- 1b8e0
		x"1d7c0001", -- 1b8e4
		x"ffff603c", -- 1b8e8
		x"206e000e", -- 1b8ec
		x"202e000a", -- 1b8f0
		x"54807200", -- 1b8f4
		x"12300800", -- 1b8f8
		x"e34148c1", -- 1b8fc
		x"2d41fffa", -- 1b900
		x"66081d7c", -- 1b904
		x"0001ffff", -- 1b908
		x"601a202e", -- 1b90c
		x"fffad1ae", -- 1b910
		x"000a0cae", -- 1b914
		x"00000fff", -- 1b918
		x"000a5ec0", -- 1b91c
		x"02000001", -- 1b920
		x"1d40ffff", -- 1b924
		x"4a2effff", -- 1b928
		x"67882d6e", -- 1b92c
		x"000a0012", -- 1b930
		x"4e5e205f", -- 1b934
		x"defc000a", -- 1b938
		x"4ed04e56", -- 1b93c
		x"fff8246e", -- 1b940
		x"001014bc", -- 1b944
		x"0000206e", -- 1b948
		x"000c4290", -- 1b94c
		x"598f2f2e", -- 1b950
		x"001a2f2e", -- 1b954
		x"00161f3c", -- 1b958
		x"00044eba", -- 1b95c
		x"e7cc2d5f", -- 1b960
		x"fffa6f72", -- 1b964
		x"598f2f2e", -- 1b968
		x"001a2f2e", -- 1b96c
		x"fffa1f2e", -- 1b970
		x"00144eba", -- 1b974
		x"ff2e206e", -- 1b978
		x"000c209f", -- 1b97c
		x"206e000c", -- 1b980
		x"4a906f52", -- 1b984
		x"206e001a", -- 1b988
		x"226e000c", -- 1b98c
		x"20115880", -- 1b990
		x"1d700800", -- 1b994
		x"fff9598f", -- 1b998
		x"2f2e001a", -- 1b99c
		x"2f2e0016", -- 1b9a0
		x"1f3c0001", -- 1b9a4
		x"4ebae782", -- 1b9a8
		x"2d5ffffa", -- 1b9ac
		x"6f28598f", -- 1b9b0
		x"2f2e001a", -- 1b9b4
		x"2f2efffa", -- 1b9b8
		x"1f2efff9", -- 1b9bc
		x"4ebafaba", -- 1b9c0
		x"2d5ffffa", -- 1b9c4
		x"6f102f2e", -- 1b9c8
		x"001a2f2e", -- 1b9cc
		x"fffa2f2e", -- 1b9d0
		x"00104eba", -- 1b9d4
		x"fb104e5e", -- 1b9d8
		x"205fdefc", -- 1b9dc
		x"00164ed0", -- 1b9e0
		x"4e56ffc2", -- 1b9e4
		x"206e0008", -- 1b9e8
		x"52a8ffee", -- 1b9ec
		x"45eeffe0", -- 1b9f0
		x"14bc0000", -- 1b9f4
		x"2f280008", -- 1b9f8
		x"2f28ffea", -- 1b9fc
		x"2268000c", -- 1ba00
		x"7010d0a8", -- 1ba04
		x"fff41f31", -- 1ba08
		x"0800486e", -- 1ba0c
		x"ffce486e", -- 1ba10
		x"ffc62f0e", -- 1ba14
		x"4ebaff24", -- 1ba18
		x"206e0008", -- 1ba1c
		x"2268000c", -- 1ba20
		x"2028fff4", -- 1ba24
		x"50807200", -- 1ba28
		x"12310800", -- 1ba2c
		x"70609240", -- 1ba30
		x"48c12d41", -- 1ba34
		x"ffca45ee", -- 1ba38
		x"ffe0204a", -- 1ba3c
		x"701a14fc", -- 1ba40
		x"002051c8", -- 1ba44
		x"fffa14bc", -- 1ba48
		x"0000226e", -- 1ba4c
		x"00082029", -- 1ba50
		x"ffee4eba", -- 1ba54
		x"de2e5688", -- 1ba58
		x"10fc0020", -- 1ba5c
		x"10fc0020", -- 1ba60
		x"43eeffce", -- 1ba64
		x"10d966fc", -- 1ba68
		x"534810bc", -- 1ba6c
		x"00204aae", -- 1ba70
		x"ffca6c16", -- 1ba74
		x"206e0008", -- 1ba78
		x"4868fffc", -- 1ba7c
		x"486effe0", -- 1ba80
		x"487afafa", -- 1ba84
		x"4ebae760", -- 1ba88
		x"605c206e", -- 1ba8c
		x"00084868", -- 1ba90
		x"fffc2f3c", -- 1ba94
		x"00000036", -- 1ba98
		x"4eb90000", -- 1ba9c
		x"0ae4206e", -- 1baa0
		x"00082d68", -- 1baa4
		x"fffcffc2", -- 1baa8
		x"226effc2", -- 1baac
		x"42a90000", -- 1bab0
		x"42290004", -- 1bab4
		x"137c0002", -- 1bab8
		x"0005137c", -- 1babc
		x"00200016", -- 1bac0
		x"136effe0", -- 1bac4
		x"0017136e", -- 1bac8
		x"ffe10018", -- 1bacc
		x"136effe2", -- 1bad0
		x"001945ee", -- 1bad4
		x"ffe047e9", -- 1bad8
		x"001a16da", -- 1badc
		x"66fc237c", -- 1bae0
		x"0001b580", -- 1bae4
		x"0006206e", -- 1bae8
		x"0008226d", -- 1baec
		x"ffe82368", -- 1baf0
		x"fffc0000", -- 1baf4
		x"2b68fffc", -- 1baf8
		x"ffe82d68", -- 1bafc
		x"fffcffc2", -- 1bb00
		x"226effc2", -- 1bb04
		x"42a9000a", -- 1bb08
		x"2368fff4", -- 1bb0c
		x"000e236e", -- 1bb10
		x"ffc60012", -- 1bb14
		x"2f28000c", -- 1bb18
		x"4868fff4", -- 1bb1c
		x"4ebae01c", -- 1bb20
		x"4e5e2e9f", -- 1bb24
		x"4e75207c", -- 1bb28
		x"00600001", -- 1bb2c
		x"7c007e00", -- 1bb30
		x"2f2dfff6", -- 1bb34
		x"487a000c", -- 1bb38
		x"2b4ffff6", -- 1bb3c
		x"4a100dc7", -- 1bb40
		x"6008487a", -- 1bb44
		x"fffe2b4f", -- 1bb48
		x"fff6d1fc", -- 1bb4c
		x"00010000", -- 1bb50
		x"52460c86", -- 1bb54
		x"0000001f", -- 1bb58
		x"66e2dffc", -- 1bb5c
		x"00000004", -- 1bb60
		x"2b47ffda", -- 1bb64
		x"2b5ffff6", -- 1bb68
		x"4e754e56", -- 1bb6c
		x"ffe62f0e", -- 1bb70
		x"4ebaffb4", -- 1bb74
		x"486dffec", -- 1bb78
		x"2f3c0000", -- 1bb7c
		x"00364eb9", -- 1bb80
		x"00000ae4", -- 1bb84
		x"2d6dffec", -- 1bb88
		x"ffe6206e", -- 1bb8c
		x"ffe642a8", -- 1bb90
		x"00004228", -- 1bb94
		x"0004117c", -- 1bb98
		x"00000005", -- 1bb9c
		x"43fa0256", -- 1bba0
		x"45e80006", -- 1bba4
		x"14d966fc", -- 1bba8
		x"224a4eba", -- 1bbac
		x"ed8c486d", -- 1bbb0
		x"ffe8487a", -- 1bbb4
		x"01864eba", -- 1bbb8
		x"e5fe206d", -- 1bbbc
		x"ffec20ad", -- 1bbc0
		x"ffe8486e", -- 1bbc4
		x"fffc487a", -- 1bbc8
		x"018c4eba", -- 1bbcc
		x"e5ea206d", -- 1bbd0
		x"ffe820ae", -- 1bbd4
		x"fffc2b6e", -- 1bbd8
		x"fffcffe8", -- 1bbdc
		x"486efffc", -- 1bbe0
		x"487a018e", -- 1bbe4
		x"4ebae5d0", -- 1bbe8
		x"206dffe8", -- 1bbec
		x"20aefffc", -- 1bbf0
		x"2b6efffc", -- 1bbf4
		x"ffe842ae", -- 1bbf8
		x"ffee598f", -- 1bbfc
		x"2f2e0008", -- 1bc00
		x"1f3c0002", -- 1bc04
		x"4ebadcea", -- 1bc08
		x"2d5fffea", -- 1bc0c
		x"598f2f2e", -- 1bc10
		x"000c1f3c", -- 1bc14
		x"00014eba", -- 1bc18
		x"dcd82d5f", -- 1bc1c
		x"fff87014", -- 1bc20
		x"d0aefff8", -- 1bc24
		x"2d40fff4", -- 1bc28
		x"422efff3", -- 1bc2c
		x"206e000c", -- 1bc30
		x"202efff4", -- 1bc34
		x"72001230", -- 1bc38
		x"08006d24", -- 1bc3c
		x"b27c0002", -- 1bc40
		x"6e1ee341", -- 1bc44
		x"303b1006", -- 1bc48
		x"4efb0002", -- 1bc4c
		x"0006000e", -- 1bc50
		x"000e1d7c", -- 1bc54
		x"0001fff3", -- 1bc58
		x"60062f0e", -- 1bc5c
		x"4ebafd82", -- 1bc60
		x"0cae0000", -- 1bc64
		x"0ffffff4", -- 1bc68
		x"6f061d7c", -- 1bc6c
		x"0001fff3", -- 1bc70
		x"4a2efff3", -- 1bc74
		x"67b6206d", -- 1bc78
		x"ffe820ae", -- 1bc7c
		x"fffc2b6e", -- 1bc80
		x"fffcffe8", -- 1bc84
		x"486efffc", -- 1bc88
		x"487a0168", -- 1bc8c
		x"4ebae528", -- 1bc90
		x"206dffe8", -- 1bc94
		x"20aefffc", -- 1bc98
		x"2b6efffc", -- 1bc9c
		x"ffe8486e", -- 1bca0
		x"fffc487a", -- 1bca4
		x"00e8487a", -- 1bca8
		x"e5964eba", -- 1bcac
		x"e53a206d", -- 1bcb0
		x"ffe820ae", -- 1bcb4
		x"fffc2b6e", -- 1bcb8
		x"fffcffe8", -- 1bcbc
		x"486efffc", -- 1bcc0
		x"487a00e0", -- 1bcc4
		x"487ae7dc", -- 1bcc8
		x"4ebae51c", -- 1bccc
		x"206dffe8", -- 1bcd0
		x"20aefffc", -- 1bcd4
		x"2b6efffc", -- 1bcd8
		x"ffe8486e", -- 1bcdc
		x"fffc487a", -- 1bce0
		x"00dc4eba", -- 1bce4
		x"e4d2206d", -- 1bce8
		x"ffe820ae", -- 1bcec
		x"fffc2b6e", -- 1bcf0
		x"fffcffe8", -- 1bcf4
		x"486efffc", -- 1bcf8
		x"487a00dd", -- 1bcfc
		x"48790001", -- 1bd00
		x"8e164eba", -- 1bd04
		x"e4e2206d", -- 1bd08
		x"ffe820ae", -- 1bd0c
		x"fffc2b6e", -- 1bd10
		x"fffcffe8", -- 1bd14
		x"486efffc", -- 1bd18
		x"487a0056", -- 1bd1c
		x"487ae872", -- 1bd20
		x"4ebae4c4", -- 1bd24
		x"206dffe8", -- 1bd28
		x"20aefffc", -- 1bd2c
		x"2b6efffc", -- 1bd30
		x"ffe84e5e", -- 1bd34
		x"205f504f", -- 1bd38
		x"4ed02020", -- 1bd3c
		x"436f6e66", -- 1bd40
		x"69677572", -- 1bd44
		x"61626c65", -- 1bd48
		x"20496e74", -- 1bd4c
		x"65726661", -- 1bd50
		x"63657300", -- 1bd54
		x"6b657973", -- 1bd58
		x"20496e74", -- 1bd5c
		x"65726661", -- 1bd60
		x"63652020", -- 1bd64
		x"53656c65", -- 1bd68
		x"63742043", -- 1bd6c
		x"6f646500", -- 1bd70
		x"2d2d2d2d", -- 1bd74
		x"2d2d2d2d", -- 1bd78
		x"2d2d2d2d", -- 1bd7c
		x"2d2d2d2d", -- 1bd80
		x"2d2d2d2d", -- 1bd84
		x"2d2d2d2d", -- 1bd88
		x"2d2d2d00", -- 1bd8c
		x"20204e20", -- 1bd90
		x"2073746f", -- 1bd94
		x"7265204e", -- 1bd98
		x"65772076", -- 1bd9c
		x"616c7565", -- 1bda0
		x"73002020", -- 1bda4
		x"44202073", -- 1bda8
		x"746f7265", -- 1bdac
		x"20446566", -- 1bdb0
		x"61756c74", -- 1bdb4
		x"2076616c", -- 1bdb8
		x"75657300", -- 1bdbc
		x"20202020", -- 1bdc0
		x"28746865", -- 1bdc4
		x"6e206379", -- 1bdc8
		x"636c6520", -- 1bdcc
		x"53505520", -- 1bdd0
		x"706f7765", -- 1bdd4
		x"72290020", -- 1bdd8
		x"20412020", -- 1bddc
		x"41626f72", -- 1bde0
		x"74207769", -- 1bde4
		x"74686f75", -- 1bde8
		x"74206368", -- 1bdec
		x"616e6765", -- 1bdf0
		x"73002000", -- 1bdf4
		x"54797065", -- 1bdf8
		x"205b6b65", -- 1bdfc
		x"795d0000", -- 1be00
		x"2f0c2878", -- 1be04
		x"fed4082c", -- 1be08
		x"0001005c", -- 1be0c
		x"6732285f", -- 1be10
		x"4e75082c", -- 1be14
		x"0004000b", -- 1be18
		x"67f60838", -- 1be1c
		x"0006feda", -- 1be20
		x"66ee082c", -- 1be24
		x"0001005c", -- 1be28
		x"67164a2c", -- 1be2c
		x"005d66e0", -- 1be30
		x"197c0001", -- 1be34
		x"005d297c", -- 1be38
		x"0001be04", -- 1be3c
		x"00c260d0", -- 1be40
		x"007c0700", -- 1be44
		x"4ff8fdac", -- 1be48
		x"08390003", -- 1be4c
		x"00400003", -- 1be50
		x"660e41fa", -- 1be54
		x"d9124eb9", -- 1be58
		x"000057cc", -- 1be5c
		x"4efafffe", -- 1be60
		x"2878fed4", -- 1be64
		x"297c0001", -- 1be68
		x"be1400c2", -- 1be6c
		x"41ec00ca", -- 1be70
		x"294800b6", -- 1be74
		x"422c00c0", -- 1be78
		x"197c0003", -- 1be7c
		x"00ba08ec", -- 1be80
		x"000000c0", -- 1be84
		x"08ec0002", -- 1be88
		x"00c008d4", -- 1be8c
		x"000408ec", -- 1be90
		x"000700c0", -- 1be94
		x"4eb90000", -- 1be98
		x"6d78027c", -- 1be9c
		x"f0ff297c", -- 1bea0
		x"fffffac0", -- 1bea4
		x"03302a6c", -- 1bea8
		x"033006ac", -- 1beac
		x"ffffffda", -- 1beb0
		x"03302e6c", -- 1beb4
		x"033004ac", -- 1beb8
		x"00002800", -- 1bebc
		x"03304eb9", -- 1bec0
		x"00004af4", -- 1bec4
		x"6160486d", -- 1bec8
		x"fff02f3c", -- 1becc
		x"00001000", -- 1bed0
		x"4eb90000", -- 1bed4
		x"0ae42f2d", -- 1bed8
		x"fff04879", -- 1bedc
		x"00408000", -- 1bee0
		x"4ebaddde", -- 1bee4
		x"42adffec", -- 1bee8
		x"42adffe8", -- 1beec
		x"2f2dfff0", -- 1bef0
		x"48790040", -- 1bef4
		x"80004eba", -- 1bef8
		x"fc723b7c", -- 1befc
		x"0001fff4", -- 1bf00
		x"1b7c0001", -- 1bf04
		x"ffe72f2d", -- 1bf08
		x"ffec1f3c", -- 1bf0c
		x"0001486d", -- 1bf10
		x"ffe74eb9", -- 1bf14
		x"000194c0", -- 1bf18
		x"4e753b7c", -- 1bf1c
		x"fff4fffe", -- 1bf20
		x"2e6dfff6", -- 1bf24
		x"4e7531fc", -- 1bf28
		x"4ef9fffa", -- 1bf2c
		x"21fc0001", -- 1bf30
		x"bf1efffc", -- 1bf34
		x"4e75ffff", -- 1bf38
		x"ffffffff", -- 1bf3c
		x"ffffffff", -- 1bf40
		x"ffffffff", -- 1bf44
		x"ffffffff", -- 1bf48
		x"ffffffff", -- 1bf4c
		x"ffffffff", -- 1bf50
		x"ffffffff", -- 1bf54
		x"ffffffff", -- 1bf58
		x"ffffffff", -- 1bf5c
		x"ffffffff", -- 1bf60
		x"ffffffff", -- 1bf64
		x"ffffffff", -- 1bf68
		x"ffffffff", -- 1bf6c
		x"ffffffff", -- 1bf70
		x"ffffffff", -- 1bf74
		x"ffffffff", -- 1bf78
		x"ffffffff", -- 1bf7c
		x"ffffffff", -- 1bf80
		x"ffffffff", -- 1bf84
		x"ffffffff", -- 1bf88
		x"ffffffff", -- 1bf8c
		x"ffffffff", -- 1bf90
		x"ffffffff", -- 1bf94
		x"ffffffff", -- 1bf98
		x"ffffffff", -- 1bf9c
		x"ffffffff", -- 1bfa0
		x"ffffffff", -- 1bfa4
		x"ffffffff", -- 1bfa8
		x"ffffffff", -- 1bfac
		x"ffffffff", -- 1bfb0
		x"ffffffff", -- 1bfb4
		x"ffffffff", -- 1bfb8
		x"ffffffff", -- 1bfbc
		x"ffffffff", -- 1bfc0
		x"ffffffff", -- 1bfc4
		x"ffffffff", -- 1bfc8
		x"ffffffff", -- 1bfcc
		x"ffffffff", -- 1bfd0
		x"ffffffff", -- 1bfd4
		x"ffffffff", -- 1bfd8
		x"ffffffff", -- 1bfdc
		x"ffffffff", -- 1bfe0
		x"ffffffff", -- 1bfe4
		x"ffffffff", -- 1bfe8
		x"ffffffff", -- 1bfec
		x"ffffffff", -- 1bff0
		x"ffffffff", -- 1bff4
		x"ffffffff", -- 1bff8
		x"0b35afad", -- 1bffc
		x"ffffffff", -- 1c000
		x"ffffffff", -- 1c004
		x"ffffffff", -- 1c008
		x"ffffffff", -- 1c00c
		x"ffffffff", -- 1c010
		x"ffffffff", -- 1c014
		x"ffffffff", -- 1c018
		x"ffffffff", -- 1c01c
		x"ffffffff", -- 1c020
		x"ffffffff", -- 1c024
		x"ffffffff", -- 1c028
		x"ffffffff", -- 1c02c
		x"ffffffff", -- 1c030
		x"ffffffff", -- 1c034
		x"ffffffff", -- 1c038
		x"ffffffff", -- 1c03c
		x"ffffffff", -- 1c040
		x"ffffffff", -- 1c044
		x"ffffffff", -- 1c048
		x"ffffffff", -- 1c04c
		x"ffffffff", -- 1c050
		x"ffffffff", -- 1c054
		x"ffffffff", -- 1c058
		x"ffffffff", -- 1c05c
		x"ffffffff", -- 1c060
		x"ffffffff", -- 1c064
		x"ffffffff", -- 1c068
		x"ffffffff", -- 1c06c
		x"ffffffff", -- 1c070
		x"ffffffff", -- 1c074
		x"ffffffff", -- 1c078
		x"ffffffff", -- 1c07c
		x"ffffffff", -- 1c080
		x"ffffffff", -- 1c084
		x"ffffffff", -- 1c088
		x"ffffffff", -- 1c08c
		x"ffffffff", -- 1c090
		x"ffffffff", -- 1c094
		x"ffffffff", -- 1c098
		x"ffffffff", -- 1c09c
		x"ffffffff", -- 1c0a0
		x"ffffffff", -- 1c0a4
		x"ffffffff", -- 1c0a8
		x"ffffffff", -- 1c0ac
		x"ffffffff", -- 1c0b0
		x"ffffffff", -- 1c0b4
		x"ffffffff", -- 1c0b8
		x"ffffffff", -- 1c0bc
		x"ffffffff", -- 1c0c0
		x"ffffffff", -- 1c0c4
		x"ffffffff", -- 1c0c8
		x"ffffffff", -- 1c0cc
		x"ffffffff", -- 1c0d0
		x"ffffffff", -- 1c0d4
		x"ffffffff", -- 1c0d8
		x"ffffffff", -- 1c0dc
		x"ffffffff", -- 1c0e0
		x"ffffffff", -- 1c0e4
		x"ffffffff", -- 1c0e8
		x"ffffffff", -- 1c0ec
		x"ffffffff", -- 1c0f0
		x"ffffffff", -- 1c0f4
		x"ffffffff", -- 1c0f8
		x"ffffffff", -- 1c0fc
		x"ffffffff", -- 1c100
		x"ffffffff", -- 1c104
		x"ffffffff", -- 1c108
		x"ffffffff", -- 1c10c
		x"ffffffff", -- 1c110
		x"ffffffff", -- 1c114
		x"ffffffff", -- 1c118
		x"ffffffff", -- 1c11c
		x"ffffffff", -- 1c120
		x"ffffffff", -- 1c124
		x"ffffffff", -- 1c128
		x"ffffffff", -- 1c12c
		x"ffffffff", -- 1c130
		x"ffffffff", -- 1c134
		x"ffffffff", -- 1c138
		x"ffffffff", -- 1c13c
		x"ffffffff", -- 1c140
		x"ffffffff", -- 1c144
		x"ffffffff", -- 1c148
		x"ffffffff", -- 1c14c
		x"ffffffff", -- 1c150
		x"ffffffff", -- 1c154
		x"ffffffff", -- 1c158
		x"ffffffff", -- 1c15c
		x"ffffffff", -- 1c160
		x"ffffffff", -- 1c164
		x"ffffffff", -- 1c168
		x"ffffffff", -- 1c16c
		x"ffffffff", -- 1c170
		x"ffffffff", -- 1c174
		x"ffffffff", -- 1c178
		x"ffffffff", -- 1c17c
		x"ffffffff", -- 1c180
		x"ffffffff", -- 1c184
		x"ffffffff", -- 1c188
		x"ffffffff", -- 1c18c
		x"ffffffff", -- 1c190
		x"ffffffff", -- 1c194
		x"ffffffff", -- 1c198
		x"ffffffff", -- 1c19c
		x"ffffffff", -- 1c1a0
		x"ffffffff", -- 1c1a4
		x"ffffffff", -- 1c1a8
		x"ffffffff", -- 1c1ac
		x"ffffffff", -- 1c1b0
		x"ffffffff", -- 1c1b4
		x"ffffffff", -- 1c1b8
		x"ffffffff", -- 1c1bc
		x"ffffffff", -- 1c1c0
		x"ffffffff", -- 1c1c4
		x"ffffffff", -- 1c1c8
		x"ffffffff", -- 1c1cc
		x"ffffffff", -- 1c1d0
		x"ffffffff", -- 1c1d4
		x"ffffffff", -- 1c1d8
		x"ffffffff", -- 1c1dc
		x"ffffffff", -- 1c1e0
		x"ffffffff", -- 1c1e4
		x"ffffffff", -- 1c1e8
		x"ffffffff", -- 1c1ec
		x"ffffffff", -- 1c1f0
		x"ffffffff", -- 1c1f4
		x"ffffffff", -- 1c1f8
		x"ffffffff", -- 1c1fc
		x"ffffffff", -- 1c200
		x"ffffffff", -- 1c204
		x"ffffffff", -- 1c208
		x"ffffffff", -- 1c20c
		x"ffffffff", -- 1c210
		x"ffffffff", -- 1c214
		x"ffffffff", -- 1c218
		x"ffffffff", -- 1c21c
		x"ffffffff", -- 1c220
		x"ffffffff", -- 1c224
		x"ffffffff", -- 1c228
		x"ffffffff", -- 1c22c
		x"ffffffff", -- 1c230
		x"ffffffff", -- 1c234
		x"ffffffff", -- 1c238
		x"ffffffff", -- 1c23c
		x"ffffffff", -- 1c240
		x"ffffffff", -- 1c244
		x"ffffffff", -- 1c248
		x"ffffffff", -- 1c24c
		x"ffffffff", -- 1c250
		x"ffffffff", -- 1c254
		x"ffffffff", -- 1c258
		x"ffffffff", -- 1c25c
		x"ffffffff", -- 1c260
		x"ffffffff", -- 1c264
		x"ffffffff", -- 1c268
		x"ffffffff", -- 1c26c
		x"ffffffff", -- 1c270
		x"ffffffff", -- 1c274
		x"ffffffff", -- 1c278
		x"ffffffff", -- 1c27c
		x"ffffffff", -- 1c280
		x"ffffffff", -- 1c284
		x"ffffffff", -- 1c288
		x"ffffffff", -- 1c28c
		x"ffffffff", -- 1c290
		x"ffffffff", -- 1c294
		x"ffffffff", -- 1c298
		x"ffffffff", -- 1c29c
		x"ffffffff", -- 1c2a0
		x"ffffffff", -- 1c2a4
		x"ffffffff", -- 1c2a8
		x"ffffffff", -- 1c2ac
		x"ffffffff", -- 1c2b0
		x"ffffffff", -- 1c2b4
		x"ffffffff", -- 1c2b8
		x"ffffffff", -- 1c2bc
		x"ffffffff", -- 1c2c0
		x"ffffffff", -- 1c2c4
		x"ffffffff", -- 1c2c8
		x"ffffffff", -- 1c2cc
		x"ffffffff", -- 1c2d0
		x"ffffffff", -- 1c2d4
		x"ffffffff", -- 1c2d8
		x"ffffffff", -- 1c2dc
		x"ffffffff", -- 1c2e0
		x"ffffffff", -- 1c2e4
		x"ffffffff", -- 1c2e8
		x"ffffffff", -- 1c2ec
		x"ffffffff", -- 1c2f0
		x"ffffffff", -- 1c2f4
		x"ffffffff", -- 1c2f8
		x"ffffffff", -- 1c2fc
		x"ffffffff", -- 1c300
		x"ffffffff", -- 1c304
		x"ffffffff", -- 1c308
		x"ffffffff", -- 1c30c
		x"ffffffff", -- 1c310
		x"ffffffff", -- 1c314
		x"ffffffff", -- 1c318
		x"ffffffff", -- 1c31c
		x"ffffffff", -- 1c320
		x"ffffffff", -- 1c324
		x"ffffffff", -- 1c328
		x"ffffffff", -- 1c32c
		x"ffffffff", -- 1c330
		x"ffffffff", -- 1c334
		x"ffffffff", -- 1c338
		x"ffffffff", -- 1c33c
		x"ffffffff", -- 1c340
		x"ffffffff", -- 1c344
		x"ffffffff", -- 1c348
		x"ffffffff", -- 1c34c
		x"ffffffff", -- 1c350
		x"ffffffff", -- 1c354
		x"ffffffff", -- 1c358
		x"ffffffff", -- 1c35c
		x"ffffffff", -- 1c360
		x"ffffffff", -- 1c364
		x"ffffffff", -- 1c368
		x"ffffffff", -- 1c36c
		x"ffffffff", -- 1c370
		x"ffffffff", -- 1c374
		x"ffffffff", -- 1c378
		x"ffffffff", -- 1c37c
		x"ffffffff", -- 1c380
		x"ffffffff", -- 1c384
		x"ffffffff", -- 1c388
		x"ffffffff", -- 1c38c
		x"ffffffff", -- 1c390
		x"ffffffff", -- 1c394
		x"ffffffff", -- 1c398
		x"ffffffff", -- 1c39c
		x"ffffffff", -- 1c3a0
		x"ffffffff", -- 1c3a4
		x"ffffffff", -- 1c3a8
		x"ffffffff", -- 1c3ac
		x"ffffffff", -- 1c3b0
		x"ffffffff", -- 1c3b4
		x"ffffffff", -- 1c3b8
		x"ffffffff", -- 1c3bc
		x"ffffffff", -- 1c3c0
		x"ffffffff", -- 1c3c4
		x"ffffffff", -- 1c3c8
		x"ffffffff", -- 1c3cc
		x"ffffffff", -- 1c3d0
		x"ffffffff", -- 1c3d4
		x"ffffffff", -- 1c3d8
		x"ffffffff", -- 1c3dc
		x"ffffffff", -- 1c3e0
		x"ffffffff", -- 1c3e4
		x"ffffffff", -- 1c3e8
		x"ffffffff", -- 1c3ec
		x"ffffffff", -- 1c3f0
		x"ffffffff", -- 1c3f4
		x"ffffffff", -- 1c3f8
		x"ffffffff", -- 1c3fc
		x"ffffffff", -- 1c400
		x"ffffffff", -- 1c404
		x"ffffffff", -- 1c408
		x"ffffffff", -- 1c40c
		x"ffffffff", -- 1c410
		x"ffffffff", -- 1c414
		x"ffffffff", -- 1c418
		x"ffffffff", -- 1c41c
		x"ffffffff", -- 1c420
		x"ffffffff", -- 1c424
		x"ffffffff", -- 1c428
		x"ffffffff", -- 1c42c
		x"ffffffff", -- 1c430
		x"ffffffff", -- 1c434
		x"ffffffff", -- 1c438
		x"ffffffff", -- 1c43c
		x"ffffffff", -- 1c440
		x"ffffffff", -- 1c444
		x"ffffffff", -- 1c448
		x"ffffffff", -- 1c44c
		x"ffffffff", -- 1c450
		x"ffffffff", -- 1c454
		x"ffffffff", -- 1c458
		x"ffffffff", -- 1c45c
		x"ffffffff", -- 1c460
		x"ffffffff", -- 1c464
		x"ffffffff", -- 1c468
		x"ffffffff", -- 1c46c
		x"ffffffff", -- 1c470
		x"ffffffff", -- 1c474
		x"ffffffff", -- 1c478
		x"ffffffff", -- 1c47c
		x"ffffffff", -- 1c480
		x"ffffffff", -- 1c484
		x"ffffffff", -- 1c488
		x"ffffffff", -- 1c48c
		x"ffffffff", -- 1c490
		x"ffffffff", -- 1c494
		x"ffffffff", -- 1c498
		x"ffffffff", -- 1c49c
		x"ffffffff", -- 1c4a0
		x"ffffffff", -- 1c4a4
		x"ffffffff", -- 1c4a8
		x"ffffffff", -- 1c4ac
		x"ffffffff", -- 1c4b0
		x"ffffffff", -- 1c4b4
		x"ffffffff", -- 1c4b8
		x"ffffffff", -- 1c4bc
		x"ffffffff", -- 1c4c0
		x"ffffffff", -- 1c4c4
		x"ffffffff", -- 1c4c8
		x"ffffffff", -- 1c4cc
		x"ffffffff", -- 1c4d0
		x"ffffffff", -- 1c4d4
		x"ffffffff", -- 1c4d8
		x"ffffffff", -- 1c4dc
		x"ffffffff", -- 1c4e0
		x"ffffffff", -- 1c4e4
		x"ffffffff", -- 1c4e8
		x"ffffffff", -- 1c4ec
		x"ffffffff", -- 1c4f0
		x"ffffffff", -- 1c4f4
		x"ffffffff", -- 1c4f8
		x"ffffffff", -- 1c4fc
		x"ffffffff", -- 1c500
		x"ffffffff", -- 1c504
		x"ffffffff", -- 1c508
		x"ffffffff", -- 1c50c
		x"ffffffff", -- 1c510
		x"ffffffff", -- 1c514
		x"ffffffff", -- 1c518
		x"ffffffff", -- 1c51c
		x"ffffffff", -- 1c520
		x"ffffffff", -- 1c524
		x"ffffffff", -- 1c528
		x"ffffffff", -- 1c52c
		x"ffffffff", -- 1c530
		x"ffffffff", -- 1c534
		x"ffffffff", -- 1c538
		x"ffffffff", -- 1c53c
		x"ffffffff", -- 1c540
		x"ffffffff", -- 1c544
		x"ffffffff", -- 1c548
		x"ffffffff", -- 1c54c
		x"ffffffff", -- 1c550
		x"ffffffff", -- 1c554
		x"ffffffff", -- 1c558
		x"ffffffff", -- 1c55c
		x"ffffffff", -- 1c560
		x"ffffffff", -- 1c564
		x"ffffffff", -- 1c568
		x"ffffffff", -- 1c56c
		x"ffffffff", -- 1c570
		x"ffffffff", -- 1c574
		x"ffffffff", -- 1c578
		x"ffffffff", -- 1c57c
		x"ffffffff", -- 1c580
		x"ffffffff", -- 1c584
		x"ffffffff", -- 1c588
		x"ffffffff", -- 1c58c
		x"ffffffff", -- 1c590
		x"ffffffff", -- 1c594
		x"ffffffff", -- 1c598
		x"ffffffff", -- 1c59c
		x"ffffffff", -- 1c5a0
		x"ffffffff", -- 1c5a4
		x"ffffffff", -- 1c5a8
		x"ffffffff", -- 1c5ac
		x"ffffffff", -- 1c5b0
		x"ffffffff", -- 1c5b4
		x"ffffffff", -- 1c5b8
		x"ffffffff", -- 1c5bc
		x"ffffffff", -- 1c5c0
		x"ffffffff", -- 1c5c4
		x"ffffffff", -- 1c5c8
		x"ffffffff", -- 1c5cc
		x"ffffffff", -- 1c5d0
		x"ffffffff", -- 1c5d4
		x"ffffffff", -- 1c5d8
		x"ffffffff", -- 1c5dc
		x"ffffffff", -- 1c5e0
		x"ffffffff", -- 1c5e4
		x"ffffffff", -- 1c5e8
		x"ffffffff", -- 1c5ec
		x"ffffffff", -- 1c5f0
		x"ffffffff", -- 1c5f4
		x"ffffffff", -- 1c5f8
		x"ffffffff", -- 1c5fc
		x"ffffffff", -- 1c600
		x"ffffffff", -- 1c604
		x"ffffffff", -- 1c608
		x"ffffffff", -- 1c60c
		x"ffffffff", -- 1c610
		x"ffffffff", -- 1c614
		x"ffffffff", -- 1c618
		x"ffffffff", -- 1c61c
		x"ffffffff", -- 1c620
		x"ffffffff", -- 1c624
		x"ffffffff", -- 1c628
		x"ffffffff", -- 1c62c
		x"ffffffff", -- 1c630
		x"ffffffff", -- 1c634
		x"ffffffff", -- 1c638
		x"ffffffff", -- 1c63c
		x"ffffffff", -- 1c640
		x"ffffffff", -- 1c644
		x"ffffffff", -- 1c648
		x"ffffffff", -- 1c64c
		x"ffffffff", -- 1c650
		x"ffffffff", -- 1c654
		x"ffffffff", -- 1c658
		x"ffffffff", -- 1c65c
		x"ffffffff", -- 1c660
		x"ffffffff", -- 1c664
		x"ffffffff", -- 1c668
		x"ffffffff", -- 1c66c
		x"ffffffff", -- 1c670
		x"ffffffff", -- 1c674
		x"ffffffff", -- 1c678
		x"ffffffff", -- 1c67c
		x"ffffffff", -- 1c680
		x"ffffffff", -- 1c684
		x"ffffffff", -- 1c688
		x"ffffffff", -- 1c68c
		x"ffffffff", -- 1c690
		x"ffffffff", -- 1c694
		x"ffffffff", -- 1c698
		x"ffffffff", -- 1c69c
		x"ffffffff", -- 1c6a0
		x"ffffffff", -- 1c6a4
		x"ffffffff", -- 1c6a8
		x"ffffffff", -- 1c6ac
		x"ffffffff", -- 1c6b0
		x"ffffffff", -- 1c6b4
		x"ffffffff", -- 1c6b8
		x"ffffffff", -- 1c6bc
		x"ffffffff", -- 1c6c0
		x"ffffffff", -- 1c6c4
		x"ffffffff", -- 1c6c8
		x"ffffffff", -- 1c6cc
		x"ffffffff", -- 1c6d0
		x"ffffffff", -- 1c6d4
		x"ffffffff", -- 1c6d8
		x"ffffffff", -- 1c6dc
		x"ffffffff", -- 1c6e0
		x"ffffffff", -- 1c6e4
		x"ffffffff", -- 1c6e8
		x"ffffffff", -- 1c6ec
		x"ffffffff", -- 1c6f0
		x"ffffffff", -- 1c6f4
		x"ffffffff", -- 1c6f8
		x"ffffffff", -- 1c6fc
		x"ffffffff", -- 1c700
		x"ffffffff", -- 1c704
		x"ffffffff", -- 1c708
		x"ffffffff", -- 1c70c
		x"ffffffff", -- 1c710
		x"ffffffff", -- 1c714
		x"ffffffff", -- 1c718
		x"ffffffff", -- 1c71c
		x"ffffffff", -- 1c720
		x"ffffffff", -- 1c724
		x"ffffffff", -- 1c728
		x"ffffffff", -- 1c72c
		x"ffffffff", -- 1c730
		x"ffffffff", -- 1c734
		x"ffffffff", -- 1c738
		x"ffffffff", -- 1c73c
		x"ffffffff", -- 1c740
		x"ffffffff", -- 1c744
		x"ffffffff", -- 1c748
		x"ffffffff", -- 1c74c
		x"ffffffff", -- 1c750
		x"ffffffff", -- 1c754
		x"ffffffff", -- 1c758
		x"ffffffff", -- 1c75c
		x"ffffffff", -- 1c760
		x"ffffffff", -- 1c764
		x"ffffffff", -- 1c768
		x"ffffffff", -- 1c76c
		x"ffffffff", -- 1c770
		x"ffffffff", -- 1c774
		x"ffffffff", -- 1c778
		x"ffffffff", -- 1c77c
		x"ffffffff", -- 1c780
		x"ffffffff", -- 1c784
		x"ffffffff", -- 1c788
		x"ffffffff", -- 1c78c
		x"ffffffff", -- 1c790
		x"ffffffff", -- 1c794
		x"ffffffff", -- 1c798
		x"ffffffff", -- 1c79c
		x"ffffffff", -- 1c7a0
		x"ffffffff", -- 1c7a4
		x"ffffffff", -- 1c7a8
		x"ffffffff", -- 1c7ac
		x"ffffffff", -- 1c7b0
		x"ffffffff", -- 1c7b4
		x"ffffffff", -- 1c7b8
		x"ffffffff", -- 1c7bc
		x"ffffffff", -- 1c7c0
		x"ffffffff", -- 1c7c4
		x"ffffffff", -- 1c7c8
		x"ffffffff", -- 1c7cc
		x"ffffffff", -- 1c7d0
		x"ffffffff", -- 1c7d4
		x"ffffffff", -- 1c7d8
		x"ffffffff", -- 1c7dc
		x"ffffffff", -- 1c7e0
		x"ffffffff", -- 1c7e4
		x"ffffffff", -- 1c7e8
		x"ffffffff", -- 1c7ec
		x"ffffffff", -- 1c7f0
		x"ffffffff", -- 1c7f4
		x"ffffffff", -- 1c7f8
		x"ffffffff", -- 1c7fc
		x"ffffffff", -- 1c800
		x"ffffffff", -- 1c804
		x"ffffffff", -- 1c808
		x"ffffffff", -- 1c80c
		x"ffffffff", -- 1c810
		x"ffffffff", -- 1c814
		x"ffffffff", -- 1c818
		x"ffffffff", -- 1c81c
		x"ffffffff", -- 1c820
		x"ffffffff", -- 1c824
		x"ffffffff", -- 1c828
		x"ffffffff", -- 1c82c
		x"ffffffff", -- 1c830
		x"ffffffff", -- 1c834
		x"ffffffff", -- 1c838
		x"ffffffff", -- 1c83c
		x"ffffffff", -- 1c840
		x"ffffffff", -- 1c844
		x"ffffffff", -- 1c848
		x"ffffffff", -- 1c84c
		x"ffffffff", -- 1c850
		x"ffffffff", -- 1c854
		x"ffffffff", -- 1c858
		x"ffffffff", -- 1c85c
		x"ffffffff", -- 1c860
		x"ffffffff", -- 1c864
		x"ffffffff", -- 1c868
		x"ffffffff", -- 1c86c
		x"ffffffff", -- 1c870
		x"ffffffff", -- 1c874
		x"ffffffff", -- 1c878
		x"ffffffff", -- 1c87c
		x"ffffffff", -- 1c880
		x"ffffffff", -- 1c884
		x"ffffffff", -- 1c888
		x"ffffffff", -- 1c88c
		x"ffffffff", -- 1c890
		x"ffffffff", -- 1c894
		x"ffffffff", -- 1c898
		x"ffffffff", -- 1c89c
		x"ffffffff", -- 1c8a0
		x"ffffffff", -- 1c8a4
		x"ffffffff", -- 1c8a8
		x"ffffffff", -- 1c8ac
		x"ffffffff", -- 1c8b0
		x"ffffffff", -- 1c8b4
		x"ffffffff", -- 1c8b8
		x"ffffffff", -- 1c8bc
		x"ffffffff", -- 1c8c0
		x"ffffffff", -- 1c8c4
		x"ffffffff", -- 1c8c8
		x"ffffffff", -- 1c8cc
		x"ffffffff", -- 1c8d0
		x"ffffffff", -- 1c8d4
		x"ffffffff", -- 1c8d8
		x"ffffffff", -- 1c8dc
		x"ffffffff", -- 1c8e0
		x"ffffffff", -- 1c8e4
		x"ffffffff", -- 1c8e8
		x"ffffffff", -- 1c8ec
		x"ffffffff", -- 1c8f0
		x"ffffffff", -- 1c8f4
		x"ffffffff", -- 1c8f8
		x"ffffffff", -- 1c8fc
		x"ffffffff", -- 1c900
		x"ffffffff", -- 1c904
		x"ffffffff", -- 1c908
		x"ffffffff", -- 1c90c
		x"ffffffff", -- 1c910
		x"ffffffff", -- 1c914
		x"ffffffff", -- 1c918
		x"ffffffff", -- 1c91c
		x"ffffffff", -- 1c920
		x"ffffffff", -- 1c924
		x"ffffffff", -- 1c928
		x"ffffffff", -- 1c92c
		x"ffffffff", -- 1c930
		x"ffffffff", -- 1c934
		x"ffffffff", -- 1c938
		x"ffffffff", -- 1c93c
		x"ffffffff", -- 1c940
		x"ffffffff", -- 1c944
		x"ffffffff", -- 1c948
		x"ffffffff", -- 1c94c
		x"ffffffff", -- 1c950
		x"ffffffff", -- 1c954
		x"ffffffff", -- 1c958
		x"ffffffff", -- 1c95c
		x"ffffffff", -- 1c960
		x"ffffffff", -- 1c964
		x"ffffffff", -- 1c968
		x"ffffffff", -- 1c96c
		x"ffffffff", -- 1c970
		x"ffffffff", -- 1c974
		x"ffffffff", -- 1c978
		x"ffffffff", -- 1c97c
		x"ffffffff", -- 1c980
		x"ffffffff", -- 1c984
		x"ffffffff", -- 1c988
		x"ffffffff", -- 1c98c
		x"ffffffff", -- 1c990
		x"ffffffff", -- 1c994
		x"ffffffff", -- 1c998
		x"ffffffff", -- 1c99c
		x"ffffffff", -- 1c9a0
		x"ffffffff", -- 1c9a4
		x"ffffffff", -- 1c9a8
		x"ffffffff", -- 1c9ac
		x"ffffffff", -- 1c9b0
		x"ffffffff", -- 1c9b4
		x"ffffffff", -- 1c9b8
		x"ffffffff", -- 1c9bc
		x"ffffffff", -- 1c9c0
		x"ffffffff", -- 1c9c4
		x"ffffffff", -- 1c9c8
		x"ffffffff", -- 1c9cc
		x"ffffffff", -- 1c9d0
		x"ffffffff", -- 1c9d4
		x"ffffffff", -- 1c9d8
		x"ffffffff", -- 1c9dc
		x"ffffffff", -- 1c9e0
		x"ffffffff", -- 1c9e4
		x"ffffffff", -- 1c9e8
		x"ffffffff", -- 1c9ec
		x"ffffffff", -- 1c9f0
		x"ffffffff", -- 1c9f4
		x"ffffffff", -- 1c9f8
		x"ffffffff", -- 1c9fc
		x"ffffffff", -- 1ca00
		x"ffffffff", -- 1ca04
		x"ffffffff", -- 1ca08
		x"ffffffff", -- 1ca0c
		x"ffffffff", -- 1ca10
		x"ffffffff", -- 1ca14
		x"ffffffff", -- 1ca18
		x"ffffffff", -- 1ca1c
		x"ffffffff", -- 1ca20
		x"ffffffff", -- 1ca24
		x"ffffffff", -- 1ca28
		x"ffffffff", -- 1ca2c
		x"ffffffff", -- 1ca30
		x"ffffffff", -- 1ca34
		x"ffffffff", -- 1ca38
		x"ffffffff", -- 1ca3c
		x"ffffffff", -- 1ca40
		x"ffffffff", -- 1ca44
		x"ffffffff", -- 1ca48
		x"ffffffff", -- 1ca4c
		x"ffffffff", -- 1ca50
		x"ffffffff", -- 1ca54
		x"ffffffff", -- 1ca58
		x"ffffffff", -- 1ca5c
		x"ffffffff", -- 1ca60
		x"ffffffff", -- 1ca64
		x"ffffffff", -- 1ca68
		x"ffffffff", -- 1ca6c
		x"ffffffff", -- 1ca70
		x"ffffffff", -- 1ca74
		x"ffffffff", -- 1ca78
		x"ffffffff", -- 1ca7c
		x"ffffffff", -- 1ca80
		x"ffffffff", -- 1ca84
		x"ffffffff", -- 1ca88
		x"ffffffff", -- 1ca8c
		x"ffffffff", -- 1ca90
		x"ffffffff", -- 1ca94
		x"ffffffff", -- 1ca98
		x"ffffffff", -- 1ca9c
		x"ffffffff", -- 1caa0
		x"ffffffff", -- 1caa4
		x"ffffffff", -- 1caa8
		x"ffffffff", -- 1caac
		x"ffffffff", -- 1cab0
		x"ffffffff", -- 1cab4
		x"ffffffff", -- 1cab8
		x"ffffffff", -- 1cabc
		x"ffffffff", -- 1cac0
		x"ffffffff", -- 1cac4
		x"ffffffff", -- 1cac8
		x"ffffffff", -- 1cacc
		x"ffffffff", -- 1cad0
		x"ffffffff", -- 1cad4
		x"ffffffff", -- 1cad8
		x"ffffffff", -- 1cadc
		x"ffffffff", -- 1cae0
		x"ffffffff", -- 1cae4
		x"ffffffff", -- 1cae8
		x"ffffffff", -- 1caec
		x"ffffffff", -- 1caf0
		x"ffffffff", -- 1caf4
		x"ffffffff", -- 1caf8
		x"ffffffff", -- 1cafc
		x"ffffffff", -- 1cb00
		x"ffffffff", -- 1cb04
		x"ffffffff", -- 1cb08
		x"ffffffff", -- 1cb0c
		x"ffffffff", -- 1cb10
		x"ffffffff", -- 1cb14
		x"ffffffff", -- 1cb18
		x"ffffffff", -- 1cb1c
		x"ffffffff", -- 1cb20
		x"ffffffff", -- 1cb24
		x"ffffffff", -- 1cb28
		x"ffffffff", -- 1cb2c
		x"ffffffff", -- 1cb30
		x"ffffffff", -- 1cb34
		x"ffffffff", -- 1cb38
		x"ffffffff", -- 1cb3c
		x"ffffffff", -- 1cb40
		x"ffffffff", -- 1cb44
		x"ffffffff", -- 1cb48
		x"ffffffff", -- 1cb4c
		x"ffffffff", -- 1cb50
		x"ffffffff", -- 1cb54
		x"ffffffff", -- 1cb58
		x"ffffffff", -- 1cb5c
		x"ffffffff", -- 1cb60
		x"ffffffff", -- 1cb64
		x"ffffffff", -- 1cb68
		x"ffffffff", -- 1cb6c
		x"ffffffff", -- 1cb70
		x"ffffffff", -- 1cb74
		x"ffffffff", -- 1cb78
		x"ffffffff", -- 1cb7c
		x"ffffffff", -- 1cb80
		x"ffffffff", -- 1cb84
		x"ffffffff", -- 1cb88
		x"ffffffff", -- 1cb8c
		x"ffffffff", -- 1cb90
		x"ffffffff", -- 1cb94
		x"ffffffff", -- 1cb98
		x"ffffffff", -- 1cb9c
		x"ffffffff", -- 1cba0
		x"ffffffff", -- 1cba4
		x"ffffffff", -- 1cba8
		x"ffffffff", -- 1cbac
		x"ffffffff", -- 1cbb0
		x"ffffffff", -- 1cbb4
		x"ffffffff", -- 1cbb8
		x"ffffffff", -- 1cbbc
		x"ffffffff", -- 1cbc0
		x"ffffffff", -- 1cbc4
		x"ffffffff", -- 1cbc8
		x"ffffffff", -- 1cbcc
		x"ffffffff", -- 1cbd0
		x"ffffffff", -- 1cbd4
		x"ffffffff", -- 1cbd8
		x"ffffffff", -- 1cbdc
		x"ffffffff", -- 1cbe0
		x"ffffffff", -- 1cbe4
		x"ffffffff", -- 1cbe8
		x"ffffffff", -- 1cbec
		x"ffffffff", -- 1cbf0
		x"ffffffff", -- 1cbf4
		x"ffffffff", -- 1cbf8
		x"ffffffff", -- 1cbfc
		x"ffffffff", -- 1cc00
		x"ffffffff", -- 1cc04
		x"ffffffff", -- 1cc08
		x"ffffffff", -- 1cc0c
		x"ffffffff", -- 1cc10
		x"ffffffff", -- 1cc14
		x"ffffffff", -- 1cc18
		x"ffffffff", -- 1cc1c
		x"ffffffff", -- 1cc20
		x"ffffffff", -- 1cc24
		x"ffffffff", -- 1cc28
		x"ffffffff", -- 1cc2c
		x"ffffffff", -- 1cc30
		x"ffffffff", -- 1cc34
		x"ffffffff", -- 1cc38
		x"ffffffff", -- 1cc3c
		x"ffffffff", -- 1cc40
		x"ffffffff", -- 1cc44
		x"ffffffff", -- 1cc48
		x"ffffffff", -- 1cc4c
		x"ffffffff", -- 1cc50
		x"ffffffff", -- 1cc54
		x"ffffffff", -- 1cc58
		x"ffffffff", -- 1cc5c
		x"ffffffff", -- 1cc60
		x"ffffffff", -- 1cc64
		x"ffffffff", -- 1cc68
		x"ffffffff", -- 1cc6c
		x"ffffffff", -- 1cc70
		x"ffffffff", -- 1cc74
		x"ffffffff", -- 1cc78
		x"ffffffff", -- 1cc7c
		x"ffffffff", -- 1cc80
		x"ffffffff", -- 1cc84
		x"ffffffff", -- 1cc88
		x"ffffffff", -- 1cc8c
		x"ffffffff", -- 1cc90
		x"ffffffff", -- 1cc94
		x"ffffffff", -- 1cc98
		x"ffffffff", -- 1cc9c
		x"ffffffff", -- 1cca0
		x"ffffffff", -- 1cca4
		x"ffffffff", -- 1cca8
		x"ffffffff", -- 1ccac
		x"ffffffff", -- 1ccb0
		x"ffffffff", -- 1ccb4
		x"ffffffff", -- 1ccb8
		x"ffffffff", -- 1ccbc
		x"ffffffff", -- 1ccc0
		x"ffffffff", -- 1ccc4
		x"ffffffff", -- 1ccc8
		x"ffffffff", -- 1cccc
		x"ffffffff", -- 1ccd0
		x"ffffffff", -- 1ccd4
		x"ffffffff", -- 1ccd8
		x"ffffffff", -- 1ccdc
		x"ffffffff", -- 1cce0
		x"ffffffff", -- 1cce4
		x"ffffffff", -- 1cce8
		x"ffffffff", -- 1ccec
		x"ffffffff", -- 1ccf0
		x"ffffffff", -- 1ccf4
		x"ffffffff", -- 1ccf8
		x"ffffffff", -- 1ccfc
		x"ffffffff", -- 1cd00
		x"ffffffff", -- 1cd04
		x"ffffffff", -- 1cd08
		x"ffffffff", -- 1cd0c
		x"ffffffff", -- 1cd10
		x"ffffffff", -- 1cd14
		x"ffffffff", -- 1cd18
		x"ffffffff", -- 1cd1c
		x"ffffffff", -- 1cd20
		x"ffffffff", -- 1cd24
		x"ffffffff", -- 1cd28
		x"ffffffff", -- 1cd2c
		x"ffffffff", -- 1cd30
		x"ffffffff", -- 1cd34
		x"ffffffff", -- 1cd38
		x"ffffffff", -- 1cd3c
		x"ffffffff", -- 1cd40
		x"ffffffff", -- 1cd44
		x"ffffffff", -- 1cd48
		x"ffffffff", -- 1cd4c
		x"ffffffff", -- 1cd50
		x"ffffffff", -- 1cd54
		x"ffffffff", -- 1cd58
		x"ffffffff", -- 1cd5c
		x"ffffffff", -- 1cd60
		x"ffffffff", -- 1cd64
		x"ffffffff", -- 1cd68
		x"ffffffff", -- 1cd6c
		x"ffffffff", -- 1cd70
		x"ffffffff", -- 1cd74
		x"ffffffff", -- 1cd78
		x"ffffffff", -- 1cd7c
		x"ffffffff", -- 1cd80
		x"ffffffff", -- 1cd84
		x"ffffffff", -- 1cd88
		x"ffffffff", -- 1cd8c
		x"ffffffff", -- 1cd90
		x"ffffffff", -- 1cd94
		x"ffffffff", -- 1cd98
		x"ffffffff", -- 1cd9c
		x"ffffffff", -- 1cda0
		x"ffffffff", -- 1cda4
		x"ffffffff", -- 1cda8
		x"ffffffff", -- 1cdac
		x"ffffffff", -- 1cdb0
		x"ffffffff", -- 1cdb4
		x"ffffffff", -- 1cdb8
		x"ffffffff", -- 1cdbc
		x"ffffffff", -- 1cdc0
		x"ffffffff", -- 1cdc4
		x"ffffffff", -- 1cdc8
		x"ffffffff", -- 1cdcc
		x"ffffffff", -- 1cdd0
		x"ffffffff", -- 1cdd4
		x"ffffffff", -- 1cdd8
		x"ffffffff", -- 1cddc
		x"ffffffff", -- 1cde0
		x"ffffffff", -- 1cde4
		x"ffffffff", -- 1cde8
		x"ffffffff", -- 1cdec
		x"ffffffff", -- 1cdf0
		x"ffffffff", -- 1cdf4
		x"ffffffff", -- 1cdf8
		x"ffffffff", -- 1cdfc
		x"ffffffff", -- 1ce00
		x"ffffffff", -- 1ce04
		x"ffffffff", -- 1ce08
		x"ffffffff", -- 1ce0c
		x"ffffffff", -- 1ce10
		x"ffffffff", -- 1ce14
		x"ffffffff", -- 1ce18
		x"ffffffff", -- 1ce1c
		x"ffffffff", -- 1ce20
		x"ffffffff", -- 1ce24
		x"ffffffff", -- 1ce28
		x"ffffffff", -- 1ce2c
		x"ffffffff", -- 1ce30
		x"ffffffff", -- 1ce34
		x"ffffffff", -- 1ce38
		x"ffffffff", -- 1ce3c
		x"ffffffff", -- 1ce40
		x"ffffffff", -- 1ce44
		x"ffffffff", -- 1ce48
		x"ffffffff", -- 1ce4c
		x"ffffffff", -- 1ce50
		x"ffffffff", -- 1ce54
		x"ffffffff", -- 1ce58
		x"ffffffff", -- 1ce5c
		x"ffffffff", -- 1ce60
		x"ffffffff", -- 1ce64
		x"ffffffff", -- 1ce68
		x"ffffffff", -- 1ce6c
		x"ffffffff", -- 1ce70
		x"ffffffff", -- 1ce74
		x"ffffffff", -- 1ce78
		x"ffffffff", -- 1ce7c
		x"ffffffff", -- 1ce80
		x"ffffffff", -- 1ce84
		x"ffffffff", -- 1ce88
		x"ffffffff", -- 1ce8c
		x"ffffffff", -- 1ce90
		x"ffffffff", -- 1ce94
		x"ffffffff", -- 1ce98
		x"ffffffff", -- 1ce9c
		x"ffffffff", -- 1cea0
		x"ffffffff", -- 1cea4
		x"ffffffff", -- 1cea8
		x"ffffffff", -- 1ceac
		x"ffffffff", -- 1ceb0
		x"ffffffff", -- 1ceb4
		x"ffffffff", -- 1ceb8
		x"ffffffff", -- 1cebc
		x"ffffffff", -- 1cec0
		x"ffffffff", -- 1cec4
		x"ffffffff", -- 1cec8
		x"ffffffff", -- 1cecc
		x"ffffffff", -- 1ced0
		x"ffffffff", -- 1ced4
		x"ffffffff", -- 1ced8
		x"ffffffff", -- 1cedc
		x"ffffffff", -- 1cee0
		x"ffffffff", -- 1cee4
		x"ffffffff", -- 1cee8
		x"ffffffff", -- 1ceec
		x"ffffffff", -- 1cef0
		x"ffffffff", -- 1cef4
		x"ffffffff", -- 1cef8
		x"ffffffff", -- 1cefc
		x"ffffffff", -- 1cf00
		x"ffffffff", -- 1cf04
		x"ffffffff", -- 1cf08
		x"ffffffff", -- 1cf0c
		x"ffffffff", -- 1cf10
		x"ffffffff", -- 1cf14
		x"ffffffff", -- 1cf18
		x"ffffffff", -- 1cf1c
		x"ffffffff", -- 1cf20
		x"ffffffff", -- 1cf24
		x"ffffffff", -- 1cf28
		x"ffffffff", -- 1cf2c
		x"ffffffff", -- 1cf30
		x"ffffffff", -- 1cf34
		x"ffffffff", -- 1cf38
		x"ffffffff", -- 1cf3c
		x"ffffffff", -- 1cf40
		x"ffffffff", -- 1cf44
		x"ffffffff", -- 1cf48
		x"ffffffff", -- 1cf4c
		x"ffffffff", -- 1cf50
		x"ffffffff", -- 1cf54
		x"ffffffff", -- 1cf58
		x"ffffffff", -- 1cf5c
		x"ffffffff", -- 1cf60
		x"ffffffff", -- 1cf64
		x"ffffffff", -- 1cf68
		x"ffffffff", -- 1cf6c
		x"ffffffff", -- 1cf70
		x"ffffffff", -- 1cf74
		x"ffffffff", -- 1cf78
		x"ffffffff", -- 1cf7c
		x"ffffffff", -- 1cf80
		x"ffffffff", -- 1cf84
		x"ffffffff", -- 1cf88
		x"ffffffff", -- 1cf8c
		x"ffffffff", -- 1cf90
		x"ffffffff", -- 1cf94
		x"ffffffff", -- 1cf98
		x"ffffffff", -- 1cf9c
		x"ffffffff", -- 1cfa0
		x"ffffffff", -- 1cfa4
		x"ffffffff", -- 1cfa8
		x"ffffffff", -- 1cfac
		x"ffffffff", -- 1cfb0
		x"ffffffff", -- 1cfb4
		x"ffffffff", -- 1cfb8
		x"ffffffff", -- 1cfbc
		x"ffffffff", -- 1cfc0
		x"ffffffff", -- 1cfc4
		x"ffffffff", -- 1cfc8
		x"ffffffff", -- 1cfcc
		x"ffffffff", -- 1cfd0
		x"ffffffff", -- 1cfd4
		x"ffffffff", -- 1cfd8
		x"ffffffff", -- 1cfdc
		x"ffffffff", -- 1cfe0
		x"ffffffff", -- 1cfe4
		x"ffffffff", -- 1cfe8
		x"ffffffff", -- 1cfec
		x"ffffffff", -- 1cff0
		x"ffffffff", -- 1cff4
		x"ffffffff", -- 1cff8
		x"ffffffff", -- 1cffc
		x"ffffffff", -- 1d000
		x"ffffffff", -- 1d004
		x"ffffffff", -- 1d008
		x"ffffffff", -- 1d00c
		x"ffffffff", -- 1d010
		x"ffffffff", -- 1d014
		x"ffffffff", -- 1d018
		x"ffffffff", -- 1d01c
		x"ffffffff", -- 1d020
		x"ffffffff", -- 1d024
		x"ffffffff", -- 1d028
		x"ffffffff", -- 1d02c
		x"ffffffff", -- 1d030
		x"ffffffff", -- 1d034
		x"ffffffff", -- 1d038
		x"ffffffff", -- 1d03c
		x"ffffffff", -- 1d040
		x"ffffffff", -- 1d044
		x"ffffffff", -- 1d048
		x"ffffffff", -- 1d04c
		x"ffffffff", -- 1d050
		x"ffffffff", -- 1d054
		x"ffffffff", -- 1d058
		x"ffffffff", -- 1d05c
		x"ffffffff", -- 1d060
		x"ffffffff", -- 1d064
		x"ffffffff", -- 1d068
		x"ffffffff", -- 1d06c
		x"ffffffff", -- 1d070
		x"ffffffff", -- 1d074
		x"ffffffff", -- 1d078
		x"ffffffff", -- 1d07c
		x"ffffffff", -- 1d080
		x"ffffffff", -- 1d084
		x"ffffffff", -- 1d088
		x"ffffffff", -- 1d08c
		x"ffffffff", -- 1d090
		x"ffffffff", -- 1d094
		x"ffffffff", -- 1d098
		x"ffffffff", -- 1d09c
		x"ffffffff", -- 1d0a0
		x"ffffffff", -- 1d0a4
		x"ffffffff", -- 1d0a8
		x"ffffffff", -- 1d0ac
		x"ffffffff", -- 1d0b0
		x"ffffffff", -- 1d0b4
		x"ffffffff", -- 1d0b8
		x"ffffffff", -- 1d0bc
		x"ffffffff", -- 1d0c0
		x"ffffffff", -- 1d0c4
		x"ffffffff", -- 1d0c8
		x"ffffffff", -- 1d0cc
		x"ffffffff", -- 1d0d0
		x"ffffffff", -- 1d0d4
		x"ffffffff", -- 1d0d8
		x"ffffffff", -- 1d0dc
		x"ffffffff", -- 1d0e0
		x"ffffffff", -- 1d0e4
		x"ffffffff", -- 1d0e8
		x"ffffffff", -- 1d0ec
		x"ffffffff", -- 1d0f0
		x"ffffffff", -- 1d0f4
		x"ffffffff", -- 1d0f8
		x"ffffffff", -- 1d0fc
		x"ffffffff", -- 1d100
		x"ffffffff", -- 1d104
		x"ffffffff", -- 1d108
		x"ffffffff", -- 1d10c
		x"ffffffff", -- 1d110
		x"ffffffff", -- 1d114
		x"ffffffff", -- 1d118
		x"ffffffff", -- 1d11c
		x"ffffffff", -- 1d120
		x"ffffffff", -- 1d124
		x"ffffffff", -- 1d128
		x"ffffffff", -- 1d12c
		x"ffffffff", -- 1d130
		x"ffffffff", -- 1d134
		x"ffffffff", -- 1d138
		x"ffffffff", -- 1d13c
		x"ffffffff", -- 1d140
		x"ffffffff", -- 1d144
		x"ffffffff", -- 1d148
		x"ffffffff", -- 1d14c
		x"ffffffff", -- 1d150
		x"ffffffff", -- 1d154
		x"ffffffff", -- 1d158
		x"ffffffff", -- 1d15c
		x"ffffffff", -- 1d160
		x"ffffffff", -- 1d164
		x"ffffffff", -- 1d168
		x"ffffffff", -- 1d16c
		x"ffffffff", -- 1d170
		x"ffffffff", -- 1d174
		x"ffffffff", -- 1d178
		x"ffffffff", -- 1d17c
		x"ffffffff", -- 1d180
		x"ffffffff", -- 1d184
		x"ffffffff", -- 1d188
		x"ffffffff", -- 1d18c
		x"ffffffff", -- 1d190
		x"ffffffff", -- 1d194
		x"ffffffff", -- 1d198
		x"ffffffff", -- 1d19c
		x"ffffffff", -- 1d1a0
		x"ffffffff", -- 1d1a4
		x"ffffffff", -- 1d1a8
		x"ffffffff", -- 1d1ac
		x"ffffffff", -- 1d1b0
		x"ffffffff", -- 1d1b4
		x"ffffffff", -- 1d1b8
		x"ffffffff", -- 1d1bc
		x"ffffffff", -- 1d1c0
		x"ffffffff", -- 1d1c4
		x"ffffffff", -- 1d1c8
		x"ffffffff", -- 1d1cc
		x"ffffffff", -- 1d1d0
		x"ffffffff", -- 1d1d4
		x"ffffffff", -- 1d1d8
		x"ffffffff", -- 1d1dc
		x"ffffffff", -- 1d1e0
		x"ffffffff", -- 1d1e4
		x"ffffffff", -- 1d1e8
		x"ffffffff", -- 1d1ec
		x"ffffffff", -- 1d1f0
		x"ffffffff", -- 1d1f4
		x"ffffffff", -- 1d1f8
		x"ffffffff", -- 1d1fc
		x"ffffffff", -- 1d200
		x"ffffffff", -- 1d204
		x"ffffffff", -- 1d208
		x"ffffffff", -- 1d20c
		x"ffffffff", -- 1d210
		x"ffffffff", -- 1d214
		x"ffffffff", -- 1d218
		x"ffffffff", -- 1d21c
		x"ffffffff", -- 1d220
		x"ffffffff", -- 1d224
		x"ffffffff", -- 1d228
		x"ffffffff", -- 1d22c
		x"ffffffff", -- 1d230
		x"ffffffff", -- 1d234
		x"ffffffff", -- 1d238
		x"ffffffff", -- 1d23c
		x"ffffffff", -- 1d240
		x"ffffffff", -- 1d244
		x"ffffffff", -- 1d248
		x"ffffffff", -- 1d24c
		x"ffffffff", -- 1d250
		x"ffffffff", -- 1d254
		x"ffffffff", -- 1d258
		x"ffffffff", -- 1d25c
		x"ffffffff", -- 1d260
		x"ffffffff", -- 1d264
		x"ffffffff", -- 1d268
		x"ffffffff", -- 1d26c
		x"ffffffff", -- 1d270
		x"ffffffff", -- 1d274
		x"ffffffff", -- 1d278
		x"ffffffff", -- 1d27c
		x"ffffffff", -- 1d280
		x"ffffffff", -- 1d284
		x"ffffffff", -- 1d288
		x"ffffffff", -- 1d28c
		x"ffffffff", -- 1d290
		x"ffffffff", -- 1d294
		x"ffffffff", -- 1d298
		x"ffffffff", -- 1d29c
		x"ffffffff", -- 1d2a0
		x"ffffffff", -- 1d2a4
		x"ffffffff", -- 1d2a8
		x"ffffffff", -- 1d2ac
		x"ffffffff", -- 1d2b0
		x"ffffffff", -- 1d2b4
		x"ffffffff", -- 1d2b8
		x"ffffffff", -- 1d2bc
		x"ffffffff", -- 1d2c0
		x"ffffffff", -- 1d2c4
		x"ffffffff", -- 1d2c8
		x"ffffffff", -- 1d2cc
		x"ffffffff", -- 1d2d0
		x"ffffffff", -- 1d2d4
		x"ffffffff", -- 1d2d8
		x"ffffffff", -- 1d2dc
		x"ffffffff", -- 1d2e0
		x"ffffffff", -- 1d2e4
		x"ffffffff", -- 1d2e8
		x"ffffffff", -- 1d2ec
		x"ffffffff", -- 1d2f0
		x"ffffffff", -- 1d2f4
		x"ffffffff", -- 1d2f8
		x"ffffffff", -- 1d2fc
		x"ffffffff", -- 1d300
		x"ffffffff", -- 1d304
		x"ffffffff", -- 1d308
		x"ffffffff", -- 1d30c
		x"ffffffff", -- 1d310
		x"ffffffff", -- 1d314
		x"ffffffff", -- 1d318
		x"ffffffff", -- 1d31c
		x"ffffffff", -- 1d320
		x"ffffffff", -- 1d324
		x"ffffffff", -- 1d328
		x"ffffffff", -- 1d32c
		x"ffffffff", -- 1d330
		x"ffffffff", -- 1d334
		x"ffffffff", -- 1d338
		x"ffffffff", -- 1d33c
		x"ffffffff", -- 1d340
		x"ffffffff", -- 1d344
		x"ffffffff", -- 1d348
		x"ffffffff", -- 1d34c
		x"ffffffff", -- 1d350
		x"ffffffff", -- 1d354
		x"ffffffff", -- 1d358
		x"ffffffff", -- 1d35c
		x"ffffffff", -- 1d360
		x"ffffffff", -- 1d364
		x"ffffffff", -- 1d368
		x"ffffffff", -- 1d36c
		x"ffffffff", -- 1d370
		x"ffffffff", -- 1d374
		x"ffffffff", -- 1d378
		x"ffffffff", -- 1d37c
		x"ffffffff", -- 1d380
		x"ffffffff", -- 1d384
		x"ffffffff", -- 1d388
		x"ffffffff", -- 1d38c
		x"ffffffff", -- 1d390
		x"ffffffff", -- 1d394
		x"ffffffff", -- 1d398
		x"ffffffff", -- 1d39c
		x"ffffffff", -- 1d3a0
		x"ffffffff", -- 1d3a4
		x"ffffffff", -- 1d3a8
		x"ffffffff", -- 1d3ac
		x"ffffffff", -- 1d3b0
		x"ffffffff", -- 1d3b4
		x"ffffffff", -- 1d3b8
		x"ffffffff", -- 1d3bc
		x"ffffffff", -- 1d3c0
		x"ffffffff", -- 1d3c4
		x"ffffffff", -- 1d3c8
		x"ffffffff", -- 1d3cc
		x"ffffffff", -- 1d3d0
		x"ffffffff", -- 1d3d4
		x"ffffffff", -- 1d3d8
		x"ffffffff", -- 1d3dc
		x"ffffffff", -- 1d3e0
		x"ffffffff", -- 1d3e4
		x"ffffffff", -- 1d3e8
		x"ffffffff", -- 1d3ec
		x"ffffffff", -- 1d3f0
		x"ffffffff", -- 1d3f4
		x"ffffffff", -- 1d3f8
		x"ffffffff", -- 1d3fc
		x"ffffffff", -- 1d400
		x"ffffffff", -- 1d404
		x"ffffffff", -- 1d408
		x"ffffffff", -- 1d40c
		x"ffffffff", -- 1d410
		x"ffffffff", -- 1d414
		x"ffffffff", -- 1d418
		x"ffffffff", -- 1d41c
		x"ffffffff", -- 1d420
		x"ffffffff", -- 1d424
		x"ffffffff", -- 1d428
		x"ffffffff", -- 1d42c
		x"ffffffff", -- 1d430
		x"ffffffff", -- 1d434
		x"ffffffff", -- 1d438
		x"ffffffff", -- 1d43c
		x"ffffffff", -- 1d440
		x"ffffffff", -- 1d444
		x"ffffffff", -- 1d448
		x"ffffffff", -- 1d44c
		x"ffffffff", -- 1d450
		x"ffffffff", -- 1d454
		x"ffffffff", -- 1d458
		x"ffffffff", -- 1d45c
		x"ffffffff", -- 1d460
		x"ffffffff", -- 1d464
		x"ffffffff", -- 1d468
		x"ffffffff", -- 1d46c
		x"ffffffff", -- 1d470
		x"ffffffff", -- 1d474
		x"ffffffff", -- 1d478
		x"ffffffff", -- 1d47c
		x"ffffffff", -- 1d480
		x"ffffffff", -- 1d484
		x"ffffffff", -- 1d488
		x"ffffffff", -- 1d48c
		x"ffffffff", -- 1d490
		x"ffffffff", -- 1d494
		x"ffffffff", -- 1d498
		x"ffffffff", -- 1d49c
		x"ffffffff", -- 1d4a0
		x"ffffffff", -- 1d4a4
		x"ffffffff", -- 1d4a8
		x"ffffffff", -- 1d4ac
		x"ffffffff", -- 1d4b0
		x"ffffffff", -- 1d4b4
		x"ffffffff", -- 1d4b8
		x"ffffffff", -- 1d4bc
		x"ffffffff", -- 1d4c0
		x"ffffffff", -- 1d4c4
		x"ffffffff", -- 1d4c8
		x"ffffffff", -- 1d4cc
		x"ffffffff", -- 1d4d0
		x"ffffffff", -- 1d4d4
		x"ffffffff", -- 1d4d8
		x"ffffffff", -- 1d4dc
		x"ffffffff", -- 1d4e0
		x"ffffffff", -- 1d4e4
		x"ffffffff", -- 1d4e8
		x"ffffffff", -- 1d4ec
		x"ffffffff", -- 1d4f0
		x"ffffffff", -- 1d4f4
		x"ffffffff", -- 1d4f8
		x"ffffffff", -- 1d4fc
		x"ffffffff", -- 1d500
		x"ffffffff", -- 1d504
		x"ffffffff", -- 1d508
		x"ffffffff", -- 1d50c
		x"ffffffff", -- 1d510
		x"ffffffff", -- 1d514
		x"ffffffff", -- 1d518
		x"ffffffff", -- 1d51c
		x"ffffffff", -- 1d520
		x"ffffffff", -- 1d524
		x"ffffffff", -- 1d528
		x"ffffffff", -- 1d52c
		x"ffffffff", -- 1d530
		x"ffffffff", -- 1d534
		x"ffffffff", -- 1d538
		x"ffffffff", -- 1d53c
		x"ffffffff", -- 1d540
		x"ffffffff", -- 1d544
		x"ffffffff", -- 1d548
		x"ffffffff", -- 1d54c
		x"ffffffff", -- 1d550
		x"ffffffff", -- 1d554
		x"ffffffff", -- 1d558
		x"ffffffff", -- 1d55c
		x"ffffffff", -- 1d560
		x"ffffffff", -- 1d564
		x"ffffffff", -- 1d568
		x"ffffffff", -- 1d56c
		x"ffffffff", -- 1d570
		x"ffffffff", -- 1d574
		x"ffffffff", -- 1d578
		x"ffffffff", -- 1d57c
		x"ffffffff", -- 1d580
		x"ffffffff", -- 1d584
		x"ffffffff", -- 1d588
		x"ffffffff", -- 1d58c
		x"ffffffff", -- 1d590
		x"ffffffff", -- 1d594
		x"ffffffff", -- 1d598
		x"ffffffff", -- 1d59c
		x"ffffffff", -- 1d5a0
		x"ffffffff", -- 1d5a4
		x"ffffffff", -- 1d5a8
		x"ffffffff", -- 1d5ac
		x"ffffffff", -- 1d5b0
		x"ffffffff", -- 1d5b4
		x"ffffffff", -- 1d5b8
		x"ffffffff", -- 1d5bc
		x"ffffffff", -- 1d5c0
		x"ffffffff", -- 1d5c4
		x"ffffffff", -- 1d5c8
		x"ffffffff", -- 1d5cc
		x"ffffffff", -- 1d5d0
		x"ffffffff", -- 1d5d4
		x"ffffffff", -- 1d5d8
		x"ffffffff", -- 1d5dc
		x"ffffffff", -- 1d5e0
		x"ffffffff", -- 1d5e4
		x"ffffffff", -- 1d5e8
		x"ffffffff", -- 1d5ec
		x"ffffffff", -- 1d5f0
		x"ffffffff", -- 1d5f4
		x"ffffffff", -- 1d5f8
		x"ffffffff", -- 1d5fc
		x"ffffffff", -- 1d600
		x"ffffffff", -- 1d604
		x"ffffffff", -- 1d608
		x"ffffffff", -- 1d60c
		x"ffffffff", -- 1d610
		x"ffffffff", -- 1d614
		x"ffffffff", -- 1d618
		x"ffffffff", -- 1d61c
		x"ffffffff", -- 1d620
		x"ffffffff", -- 1d624
		x"ffffffff", -- 1d628
		x"ffffffff", -- 1d62c
		x"ffffffff", -- 1d630
		x"ffffffff", -- 1d634
		x"ffffffff", -- 1d638
		x"ffffffff", -- 1d63c
		x"ffffffff", -- 1d640
		x"ffffffff", -- 1d644
		x"ffffffff", -- 1d648
		x"ffffffff", -- 1d64c
		x"ffffffff", -- 1d650
		x"ffffffff", -- 1d654
		x"ffffffff", -- 1d658
		x"ffffffff", -- 1d65c
		x"ffffffff", -- 1d660
		x"ffffffff", -- 1d664
		x"ffffffff", -- 1d668
		x"ffffffff", -- 1d66c
		x"ffffffff", -- 1d670
		x"ffffffff", -- 1d674
		x"ffffffff", -- 1d678
		x"ffffffff", -- 1d67c
		x"ffffffff", -- 1d680
		x"ffffffff", -- 1d684
		x"ffffffff", -- 1d688
		x"ffffffff", -- 1d68c
		x"ffffffff", -- 1d690
		x"ffffffff", -- 1d694
		x"ffffffff", -- 1d698
		x"ffffffff", -- 1d69c
		x"ffffffff", -- 1d6a0
		x"ffffffff", -- 1d6a4
		x"ffffffff", -- 1d6a8
		x"ffffffff", -- 1d6ac
		x"ffffffff", -- 1d6b0
		x"ffffffff", -- 1d6b4
		x"ffffffff", -- 1d6b8
		x"ffffffff", -- 1d6bc
		x"ffffffff", -- 1d6c0
		x"ffffffff", -- 1d6c4
		x"ffffffff", -- 1d6c8
		x"ffffffff", -- 1d6cc
		x"ffffffff", -- 1d6d0
		x"ffffffff", -- 1d6d4
		x"ffffffff", -- 1d6d8
		x"ffffffff", -- 1d6dc
		x"ffffffff", -- 1d6e0
		x"ffffffff", -- 1d6e4
		x"ffffffff", -- 1d6e8
		x"ffffffff", -- 1d6ec
		x"ffffffff", -- 1d6f0
		x"ffffffff", -- 1d6f4
		x"ffffffff", -- 1d6f8
		x"ffffffff", -- 1d6fc
		x"ffffffff", -- 1d700
		x"ffffffff", -- 1d704
		x"ffffffff", -- 1d708
		x"ffffffff", -- 1d70c
		x"ffffffff", -- 1d710
		x"ffffffff", -- 1d714
		x"ffffffff", -- 1d718
		x"ffffffff", -- 1d71c
		x"ffffffff", -- 1d720
		x"ffffffff", -- 1d724
		x"ffffffff", -- 1d728
		x"ffffffff", -- 1d72c
		x"ffffffff", -- 1d730
		x"ffffffff", -- 1d734
		x"ffffffff", -- 1d738
		x"ffffffff", -- 1d73c
		x"ffffffff", -- 1d740
		x"ffffffff", -- 1d744
		x"ffffffff", -- 1d748
		x"ffffffff", -- 1d74c
		x"ffffffff", -- 1d750
		x"ffffffff", -- 1d754
		x"ffffffff", -- 1d758
		x"ffffffff", -- 1d75c
		x"ffffffff", -- 1d760
		x"ffffffff", -- 1d764
		x"ffffffff", -- 1d768
		x"ffffffff", -- 1d76c
		x"ffffffff", -- 1d770
		x"ffffffff", -- 1d774
		x"ffffffff", -- 1d778
		x"ffffffff", -- 1d77c
		x"ffffffff", -- 1d780
		x"ffffffff", -- 1d784
		x"ffffffff", -- 1d788
		x"ffffffff", -- 1d78c
		x"ffffffff", -- 1d790
		x"ffffffff", -- 1d794
		x"ffffffff", -- 1d798
		x"ffffffff", -- 1d79c
		x"ffffffff", -- 1d7a0
		x"ffffffff", -- 1d7a4
		x"ffffffff", -- 1d7a8
		x"ffffffff", -- 1d7ac
		x"ffffffff", -- 1d7b0
		x"ffffffff", -- 1d7b4
		x"ffffffff", -- 1d7b8
		x"ffffffff", -- 1d7bc
		x"ffffffff", -- 1d7c0
		x"ffffffff", -- 1d7c4
		x"ffffffff", -- 1d7c8
		x"ffffffff", -- 1d7cc
		x"ffffffff", -- 1d7d0
		x"ffffffff", -- 1d7d4
		x"ffffffff", -- 1d7d8
		x"ffffffff", -- 1d7dc
		x"ffffffff", -- 1d7e0
		x"ffffffff", -- 1d7e4
		x"ffffffff", -- 1d7e8
		x"ffffffff", -- 1d7ec
		x"ffffffff", -- 1d7f0
		x"ffffffff", -- 1d7f4
		x"ffffffff", -- 1d7f8
		x"ffffffff", -- 1d7fc
		x"ffffffff", -- 1d800
		x"ffffffff", -- 1d804
		x"ffffffff", -- 1d808
		x"ffffffff", -- 1d80c
		x"ffffffff", -- 1d810
		x"ffffffff", -- 1d814
		x"ffffffff", -- 1d818
		x"ffffffff", -- 1d81c
		x"ffffffff", -- 1d820
		x"ffffffff", -- 1d824
		x"ffffffff", -- 1d828
		x"ffffffff", -- 1d82c
		x"ffffffff", -- 1d830
		x"ffffffff", -- 1d834
		x"ffffffff", -- 1d838
		x"ffffffff", -- 1d83c
		x"ffffffff", -- 1d840
		x"ffffffff", -- 1d844
		x"ffffffff", -- 1d848
		x"ffffffff", -- 1d84c
		x"ffffffff", -- 1d850
		x"ffffffff", -- 1d854
		x"ffffffff", -- 1d858
		x"ffffffff", -- 1d85c
		x"ffffffff", -- 1d860
		x"ffffffff", -- 1d864
		x"ffffffff", -- 1d868
		x"ffffffff", -- 1d86c
		x"ffffffff", -- 1d870
		x"ffffffff", -- 1d874
		x"ffffffff", -- 1d878
		x"ffffffff", -- 1d87c
		x"ffffffff", -- 1d880
		x"ffffffff", -- 1d884
		x"ffffffff", -- 1d888
		x"ffffffff", -- 1d88c
		x"ffffffff", -- 1d890
		x"ffffffff", -- 1d894
		x"ffffffff", -- 1d898
		x"ffffffff", -- 1d89c
		x"ffffffff", -- 1d8a0
		x"ffffffff", -- 1d8a4
		x"ffffffff", -- 1d8a8
		x"ffffffff", -- 1d8ac
		x"ffffffff", -- 1d8b0
		x"ffffffff", -- 1d8b4
		x"ffffffff", -- 1d8b8
		x"ffffffff", -- 1d8bc
		x"ffffffff", -- 1d8c0
		x"ffffffff", -- 1d8c4
		x"ffffffff", -- 1d8c8
		x"ffffffff", -- 1d8cc
		x"ffffffff", -- 1d8d0
		x"ffffffff", -- 1d8d4
		x"ffffffff", -- 1d8d8
		x"ffffffff", -- 1d8dc
		x"ffffffff", -- 1d8e0
		x"ffffffff", -- 1d8e4
		x"ffffffff", -- 1d8e8
		x"ffffffff", -- 1d8ec
		x"ffffffff", -- 1d8f0
		x"ffffffff", -- 1d8f4
		x"ffffffff", -- 1d8f8
		x"ffffffff", -- 1d8fc
		x"ffffffff", -- 1d900
		x"ffffffff", -- 1d904
		x"ffffffff", -- 1d908
		x"ffffffff", -- 1d90c
		x"ffffffff", -- 1d910
		x"ffffffff", -- 1d914
		x"ffffffff", -- 1d918
		x"ffffffff", -- 1d91c
		x"ffffffff", -- 1d920
		x"ffffffff", -- 1d924
		x"ffffffff", -- 1d928
		x"ffffffff", -- 1d92c
		x"ffffffff", -- 1d930
		x"ffffffff", -- 1d934
		x"ffffffff", -- 1d938
		x"ffffffff", -- 1d93c
		x"ffffffff", -- 1d940
		x"ffffffff", -- 1d944
		x"ffffffff", -- 1d948
		x"ffffffff", -- 1d94c
		x"ffffffff", -- 1d950
		x"ffffffff", -- 1d954
		x"ffffffff", -- 1d958
		x"ffffffff", -- 1d95c
		x"ffffffff", -- 1d960
		x"ffffffff", -- 1d964
		x"ffffffff", -- 1d968
		x"ffffffff", -- 1d96c
		x"ffffffff", -- 1d970
		x"ffffffff", -- 1d974
		x"ffffffff", -- 1d978
		x"ffffffff", -- 1d97c
		x"ffffffff", -- 1d980
		x"ffffffff", -- 1d984
		x"ffffffff", -- 1d988
		x"ffffffff", -- 1d98c
		x"ffffffff", -- 1d990
		x"ffffffff", -- 1d994
		x"ffffffff", -- 1d998
		x"ffffffff", -- 1d99c
		x"ffffffff", -- 1d9a0
		x"ffffffff", -- 1d9a4
		x"ffffffff", -- 1d9a8
		x"ffffffff", -- 1d9ac
		x"ffffffff", -- 1d9b0
		x"ffffffff", -- 1d9b4
		x"ffffffff", -- 1d9b8
		x"ffffffff", -- 1d9bc
		x"ffffffff", -- 1d9c0
		x"ffffffff", -- 1d9c4
		x"ffffffff", -- 1d9c8
		x"ffffffff", -- 1d9cc
		x"ffffffff", -- 1d9d0
		x"ffffffff", -- 1d9d4
		x"ffffffff", -- 1d9d8
		x"ffffffff", -- 1d9dc
		x"ffffffff", -- 1d9e0
		x"ffffffff", -- 1d9e4
		x"ffffffff", -- 1d9e8
		x"ffffffff", -- 1d9ec
		x"ffffffff", -- 1d9f0
		x"ffffffff", -- 1d9f4
		x"ffffffff", -- 1d9f8
		x"ffffffff", -- 1d9fc
		x"ffffffff", -- 1da00
		x"ffffffff", -- 1da04
		x"ffffffff", -- 1da08
		x"ffffffff", -- 1da0c
		x"ffffffff", -- 1da10
		x"ffffffff", -- 1da14
		x"ffffffff", -- 1da18
		x"ffffffff", -- 1da1c
		x"ffffffff", -- 1da20
		x"ffffffff", -- 1da24
		x"ffffffff", -- 1da28
		x"ffffffff", -- 1da2c
		x"ffffffff", -- 1da30
		x"ffffffff", -- 1da34
		x"ffffffff", -- 1da38
		x"ffffffff", -- 1da3c
		x"ffffffff", -- 1da40
		x"ffffffff", -- 1da44
		x"ffffffff", -- 1da48
		x"ffffffff", -- 1da4c
		x"ffffffff", -- 1da50
		x"ffffffff", -- 1da54
		x"ffffffff", -- 1da58
		x"ffffffff", -- 1da5c
		x"ffffffff", -- 1da60
		x"ffffffff", -- 1da64
		x"ffffffff", -- 1da68
		x"ffffffff", -- 1da6c
		x"ffffffff", -- 1da70
		x"ffffffff", -- 1da74
		x"ffffffff", -- 1da78
		x"ffffffff", -- 1da7c
		x"ffffffff", -- 1da80
		x"ffffffff", -- 1da84
		x"ffffffff", -- 1da88
		x"ffffffff", -- 1da8c
		x"ffffffff", -- 1da90
		x"ffffffff", -- 1da94
		x"ffffffff", -- 1da98
		x"ffffffff", -- 1da9c
		x"ffffffff", -- 1daa0
		x"ffffffff", -- 1daa4
		x"ffffffff", -- 1daa8
		x"ffffffff", -- 1daac
		x"ffffffff", -- 1dab0
		x"ffffffff", -- 1dab4
		x"ffffffff", -- 1dab8
		x"ffffffff", -- 1dabc
		x"ffffffff", -- 1dac0
		x"ffffffff", -- 1dac4
		x"ffffffff", -- 1dac8
		x"ffffffff", -- 1dacc
		x"ffffffff", -- 1dad0
		x"ffffffff", -- 1dad4
		x"ffffffff", -- 1dad8
		x"ffffffff", -- 1dadc
		x"ffffffff", -- 1dae0
		x"ffffffff", -- 1dae4
		x"ffffffff", -- 1dae8
		x"ffffffff", -- 1daec
		x"ffffffff", -- 1daf0
		x"ffffffff", -- 1daf4
		x"ffffffff", -- 1daf8
		x"ffffffff", -- 1dafc
		x"ffffffff", -- 1db00
		x"ffffffff", -- 1db04
		x"ffffffff", -- 1db08
		x"ffffffff", -- 1db0c
		x"ffffffff", -- 1db10
		x"ffffffff", -- 1db14
		x"ffffffff", -- 1db18
		x"ffffffff", -- 1db1c
		x"ffffffff", -- 1db20
		x"ffffffff", -- 1db24
		x"ffffffff", -- 1db28
		x"ffffffff", -- 1db2c
		x"ffffffff", -- 1db30
		x"ffffffff", -- 1db34
		x"ffffffff", -- 1db38
		x"ffffffff", -- 1db3c
		x"ffffffff", -- 1db40
		x"ffffffff", -- 1db44
		x"ffffffff", -- 1db48
		x"ffffffff", -- 1db4c
		x"ffffffff", -- 1db50
		x"ffffffff", -- 1db54
		x"ffffffff", -- 1db58
		x"ffffffff", -- 1db5c
		x"ffffffff", -- 1db60
		x"ffffffff", -- 1db64
		x"ffffffff", -- 1db68
		x"ffffffff", -- 1db6c
		x"ffffffff", -- 1db70
		x"ffffffff", -- 1db74
		x"ffffffff", -- 1db78
		x"ffffffff", -- 1db7c
		x"ffffffff", -- 1db80
		x"ffffffff", -- 1db84
		x"ffffffff", -- 1db88
		x"ffffffff", -- 1db8c
		x"ffffffff", -- 1db90
		x"ffffffff", -- 1db94
		x"ffffffff", -- 1db98
		x"ffffffff", -- 1db9c
		x"ffffffff", -- 1dba0
		x"ffffffff", -- 1dba4
		x"ffffffff", -- 1dba8
		x"ffffffff", -- 1dbac
		x"ffffffff", -- 1dbb0
		x"ffffffff", -- 1dbb4
		x"ffffffff", -- 1dbb8
		x"ffffffff", -- 1dbbc
		x"ffffffff", -- 1dbc0
		x"ffffffff", -- 1dbc4
		x"ffffffff", -- 1dbc8
		x"ffffffff", -- 1dbcc
		x"ffffffff", -- 1dbd0
		x"ffffffff", -- 1dbd4
		x"ffffffff", -- 1dbd8
		x"ffffffff", -- 1dbdc
		x"ffffffff", -- 1dbe0
		x"ffffffff", -- 1dbe4
		x"ffffffff", -- 1dbe8
		x"ffffffff", -- 1dbec
		x"ffffffff", -- 1dbf0
		x"ffffffff", -- 1dbf4
		x"ffffffff", -- 1dbf8
		x"ffffffff", -- 1dbfc
		x"ffffffff", -- 1dc00
		x"ffffffff", -- 1dc04
		x"ffffffff", -- 1dc08
		x"ffffffff", -- 1dc0c
		x"ffffffff", -- 1dc10
		x"ffffffff", -- 1dc14
		x"ffffffff", -- 1dc18
		x"ffffffff", -- 1dc1c
		x"ffffffff", -- 1dc20
		x"ffffffff", -- 1dc24
		x"ffffffff", -- 1dc28
		x"ffffffff", -- 1dc2c
		x"ffffffff", -- 1dc30
		x"ffffffff", -- 1dc34
		x"ffffffff", -- 1dc38
		x"ffffffff", -- 1dc3c
		x"ffffffff", -- 1dc40
		x"ffffffff", -- 1dc44
		x"ffffffff", -- 1dc48
		x"ffffffff", -- 1dc4c
		x"ffffffff", -- 1dc50
		x"ffffffff", -- 1dc54
		x"ffffffff", -- 1dc58
		x"ffffffff", -- 1dc5c
		x"ffffffff", -- 1dc60
		x"ffffffff", -- 1dc64
		x"ffffffff", -- 1dc68
		x"ffffffff", -- 1dc6c
		x"ffffffff", -- 1dc70
		x"ffffffff", -- 1dc74
		x"ffffffff", -- 1dc78
		x"ffffffff", -- 1dc7c
		x"ffffffff", -- 1dc80
		x"ffffffff", -- 1dc84
		x"ffffffff", -- 1dc88
		x"ffffffff", -- 1dc8c
		x"ffffffff", -- 1dc90
		x"ffffffff", -- 1dc94
		x"ffffffff", -- 1dc98
		x"ffffffff", -- 1dc9c
		x"ffffffff", -- 1dca0
		x"ffffffff", -- 1dca4
		x"ffffffff", -- 1dca8
		x"ffffffff", -- 1dcac
		x"ffffffff", -- 1dcb0
		x"ffffffff", -- 1dcb4
		x"ffffffff", -- 1dcb8
		x"ffffffff", -- 1dcbc
		x"ffffffff", -- 1dcc0
		x"ffffffff", -- 1dcc4
		x"ffffffff", -- 1dcc8
		x"ffffffff", -- 1dccc
		x"ffffffff", -- 1dcd0
		x"ffffffff", -- 1dcd4
		x"ffffffff", -- 1dcd8
		x"ffffffff", -- 1dcdc
		x"ffffffff", -- 1dce0
		x"ffffffff", -- 1dce4
		x"ffffffff", -- 1dce8
		x"ffffffff", -- 1dcec
		x"ffffffff", -- 1dcf0
		x"ffffffff", -- 1dcf4
		x"ffffffff", -- 1dcf8
		x"ffffffff", -- 1dcfc
		x"ffffffff", -- 1dd00
		x"ffffffff", -- 1dd04
		x"ffffffff", -- 1dd08
		x"ffffffff", -- 1dd0c
		x"ffffffff", -- 1dd10
		x"ffffffff", -- 1dd14
		x"ffffffff", -- 1dd18
		x"ffffffff", -- 1dd1c
		x"ffffffff", -- 1dd20
		x"ffffffff", -- 1dd24
		x"ffffffff", -- 1dd28
		x"ffffffff", -- 1dd2c
		x"ffffffff", -- 1dd30
		x"ffffffff", -- 1dd34
		x"ffffffff", -- 1dd38
		x"ffffffff", -- 1dd3c
		x"ffffffff", -- 1dd40
		x"ffffffff", -- 1dd44
		x"ffffffff", -- 1dd48
		x"ffffffff", -- 1dd4c
		x"ffffffff", -- 1dd50
		x"ffffffff", -- 1dd54
		x"ffffffff", -- 1dd58
		x"ffffffff", -- 1dd5c
		x"ffffffff", -- 1dd60
		x"ffffffff", -- 1dd64
		x"ffffffff", -- 1dd68
		x"ffffffff", -- 1dd6c
		x"ffffffff", -- 1dd70
		x"ffffffff", -- 1dd74
		x"ffffffff", -- 1dd78
		x"ffffffff", -- 1dd7c
		x"ffffffff", -- 1dd80
		x"ffffffff", -- 1dd84
		x"ffffffff", -- 1dd88
		x"ffffffff", -- 1dd8c
		x"ffffffff", -- 1dd90
		x"ffffffff", -- 1dd94
		x"ffffffff", -- 1dd98
		x"ffffffff", -- 1dd9c
		x"ffffffff", -- 1dda0
		x"ffffffff", -- 1dda4
		x"ffffffff", -- 1dda8
		x"ffffffff", -- 1ddac
		x"ffffffff", -- 1ddb0
		x"ffffffff", -- 1ddb4
		x"ffffffff", -- 1ddb8
		x"ffffffff", -- 1ddbc
		x"ffffffff", -- 1ddc0
		x"ffffffff", -- 1ddc4
		x"ffffffff", -- 1ddc8
		x"ffffffff", -- 1ddcc
		x"ffffffff", -- 1ddd0
		x"ffffffff", -- 1ddd4
		x"ffffffff", -- 1ddd8
		x"ffffffff", -- 1dddc
		x"ffffffff", -- 1dde0
		x"ffffffff", -- 1dde4
		x"ffffffff", -- 1dde8
		x"ffffffff", -- 1ddec
		x"ffffffff", -- 1ddf0
		x"ffffffff", -- 1ddf4
		x"ffffffff", -- 1ddf8
		x"ffffffff", -- 1ddfc
		x"ffffffff", -- 1de00
		x"ffffffff", -- 1de04
		x"ffffffff", -- 1de08
		x"ffffffff", -- 1de0c
		x"ffffffff", -- 1de10
		x"ffffffff", -- 1de14
		x"ffffffff", -- 1de18
		x"ffffffff", -- 1de1c
		x"ffffffff", -- 1de20
		x"ffffffff", -- 1de24
		x"ffffffff", -- 1de28
		x"ffffffff", -- 1de2c
		x"ffffffff", -- 1de30
		x"ffffffff", -- 1de34
		x"ffffffff", -- 1de38
		x"ffffffff", -- 1de3c
		x"ffffffff", -- 1de40
		x"ffffffff", -- 1de44
		x"ffffffff", -- 1de48
		x"ffffffff", -- 1de4c
		x"ffffffff", -- 1de50
		x"ffffffff", -- 1de54
		x"ffffffff", -- 1de58
		x"ffffffff", -- 1de5c
		x"ffffffff", -- 1de60
		x"ffffffff", -- 1de64
		x"ffffffff", -- 1de68
		x"ffffffff", -- 1de6c
		x"ffffffff", -- 1de70
		x"ffffffff", -- 1de74
		x"ffffffff", -- 1de78
		x"ffffffff", -- 1de7c
		x"ffffffff", -- 1de80
		x"ffffffff", -- 1de84
		x"ffffffff", -- 1de88
		x"ffffffff", -- 1de8c
		x"ffffffff", -- 1de90
		x"ffffffff", -- 1de94
		x"ffffffff", -- 1de98
		x"ffffffff", -- 1de9c
		x"ffffffff", -- 1dea0
		x"ffffffff", -- 1dea4
		x"ffffffff", -- 1dea8
		x"ffffffff", -- 1deac
		x"ffffffff", -- 1deb0
		x"ffffffff", -- 1deb4
		x"ffffffff", -- 1deb8
		x"ffffffff", -- 1debc
		x"ffffffff", -- 1dec0
		x"ffffffff", -- 1dec4
		x"ffffffff", -- 1dec8
		x"ffffffff", -- 1decc
		x"ffffffff", -- 1ded0
		x"ffffffff", -- 1ded4
		x"ffffffff", -- 1ded8
		x"ffffffff", -- 1dedc
		x"ffffffff", -- 1dee0
		x"ffffffff", -- 1dee4
		x"ffffffff", -- 1dee8
		x"ffffffff", -- 1deec
		x"ffffffff", -- 1def0
		x"ffffffff", -- 1def4
		x"ffffffff", -- 1def8
		x"ffffffff", -- 1defc
		x"ffffffff", -- 1df00
		x"ffffffff", -- 1df04
		x"ffffffff", -- 1df08
		x"ffffffff", -- 1df0c
		x"ffffffff", -- 1df10
		x"ffffffff", -- 1df14
		x"ffffffff", -- 1df18
		x"ffffffff", -- 1df1c
		x"ffffffff", -- 1df20
		x"ffffffff", -- 1df24
		x"ffffffff", -- 1df28
		x"ffffffff", -- 1df2c
		x"ffffffff", -- 1df30
		x"ffffffff", -- 1df34
		x"ffffffff", -- 1df38
		x"ffffffff", -- 1df3c
		x"ffffffff", -- 1df40
		x"ffffffff", -- 1df44
		x"ffffffff", -- 1df48
		x"ffffffff", -- 1df4c
		x"ffffffff", -- 1df50
		x"ffffffff", -- 1df54
		x"ffffffff", -- 1df58
		x"ffffffff", -- 1df5c
		x"ffffffff", -- 1df60
		x"ffffffff", -- 1df64
		x"ffffffff", -- 1df68
		x"ffffffff", -- 1df6c
		x"ffffffff", -- 1df70
		x"ffffffff", -- 1df74
		x"ffffffff", -- 1df78
		x"ffffffff", -- 1df7c
		x"ffffffff", -- 1df80
		x"ffffffff", -- 1df84
		x"ffffffff", -- 1df88
		x"ffffffff", -- 1df8c
		x"ffffffff", -- 1df90
		x"ffffffff", -- 1df94
		x"ffffffff", -- 1df98
		x"ffffffff", -- 1df9c
		x"ffffffff", -- 1dfa0
		x"ffffffff", -- 1dfa4
		x"ffffffff", -- 1dfa8
		x"ffffffff", -- 1dfac
		x"ffffffff", -- 1dfb0
		x"ffffffff", -- 1dfb4
		x"ffffffff", -- 1dfb8
		x"ffffffff", -- 1dfbc
		x"ffffffff", -- 1dfc0
		x"ffffffff", -- 1dfc4
		x"ffffffff", -- 1dfc8
		x"ffffffff", -- 1dfcc
		x"ffffffff", -- 1dfd0
		x"ffffffff", -- 1dfd4
		x"ffffffff", -- 1dfd8
		x"ffffffff", -- 1dfdc
		x"ffffffff", -- 1dfe0
		x"ffffffff", -- 1dfe4
		x"ffffffff", -- 1dfe8
		x"ffffffff", -- 1dfec
		x"ffffffff", -- 1dff0
		x"ffffffff", -- 1dff4
		x"ffffffff", -- 1dff8
		x"ffffffff", -- 1dffc
		x"ffffffff", -- 1e000
		x"ffffffff", -- 1e004
		x"ffffffff", -- 1e008
		x"ffffffff", -- 1e00c
		x"ffffffff", -- 1e010
		x"ffffffff", -- 1e014
		x"ffffffff", -- 1e018
		x"ffffffff", -- 1e01c
		x"ffffffff", -- 1e020
		x"ffffffff", -- 1e024
		x"ffffffff", -- 1e028
		x"ffffffff", -- 1e02c
		x"ffffffff", -- 1e030
		x"ffffffff", -- 1e034
		x"ffffffff", -- 1e038
		x"ffffffff", -- 1e03c
		x"ffffffff", -- 1e040
		x"ffffffff", -- 1e044
		x"ffffffff", -- 1e048
		x"ffffffff", -- 1e04c
		x"ffffffff", -- 1e050
		x"ffffffff", -- 1e054
		x"ffffffff", -- 1e058
		x"ffffffff", -- 1e05c
		x"ffffffff", -- 1e060
		x"ffffffff", -- 1e064
		x"ffffffff", -- 1e068
		x"ffffffff", -- 1e06c
		x"ffffffff", -- 1e070
		x"ffffffff", -- 1e074
		x"ffffffff", -- 1e078
		x"ffffffff", -- 1e07c
		x"ffffffff", -- 1e080
		x"ffffffff", -- 1e084
		x"ffffffff", -- 1e088
		x"ffffffff", -- 1e08c
		x"ffffffff", -- 1e090
		x"ffffffff", -- 1e094
		x"ffffffff", -- 1e098
		x"ffffffff", -- 1e09c
		x"ffffffff", -- 1e0a0
		x"ffffffff", -- 1e0a4
		x"ffffffff", -- 1e0a8
		x"ffffffff", -- 1e0ac
		x"ffffffff", -- 1e0b0
		x"ffffffff", -- 1e0b4
		x"ffffffff", -- 1e0b8
		x"ffffffff", -- 1e0bc
		x"ffffffff", -- 1e0c0
		x"ffffffff", -- 1e0c4
		x"ffffffff", -- 1e0c8
		x"ffffffff", -- 1e0cc
		x"ffffffff", -- 1e0d0
		x"ffffffff", -- 1e0d4
		x"ffffffff", -- 1e0d8
		x"ffffffff", -- 1e0dc
		x"ffffffff", -- 1e0e0
		x"ffffffff", -- 1e0e4
		x"ffffffff", -- 1e0e8
		x"ffffffff", -- 1e0ec
		x"ffffffff", -- 1e0f0
		x"ffffffff", -- 1e0f4
		x"ffffffff", -- 1e0f8
		x"ffffffff", -- 1e0fc
		x"ffffffff", -- 1e100
		x"ffffffff", -- 1e104
		x"ffffffff", -- 1e108
		x"ffffffff", -- 1e10c
		x"ffffffff", -- 1e110
		x"ffffffff", -- 1e114
		x"ffffffff", -- 1e118
		x"ffffffff", -- 1e11c
		x"ffffffff", -- 1e120
		x"ffffffff", -- 1e124
		x"ffffffff", -- 1e128
		x"ffffffff", -- 1e12c
		x"ffffffff", -- 1e130
		x"ffffffff", -- 1e134
		x"ffffffff", -- 1e138
		x"ffffffff", -- 1e13c
		x"ffffffff", -- 1e140
		x"ffffffff", -- 1e144
		x"ffffffff", -- 1e148
		x"ffffffff", -- 1e14c
		x"ffffffff", -- 1e150
		x"ffffffff", -- 1e154
		x"ffffffff", -- 1e158
		x"ffffffff", -- 1e15c
		x"ffffffff", -- 1e160
		x"ffffffff", -- 1e164
		x"ffffffff", -- 1e168
		x"ffffffff", -- 1e16c
		x"ffffffff", -- 1e170
		x"ffffffff", -- 1e174
		x"ffffffff", -- 1e178
		x"ffffffff", -- 1e17c
		x"ffffffff", -- 1e180
		x"ffffffff", -- 1e184
		x"ffffffff", -- 1e188
		x"ffffffff", -- 1e18c
		x"ffffffff", -- 1e190
		x"ffffffff", -- 1e194
		x"ffffffff", -- 1e198
		x"ffffffff", -- 1e19c
		x"ffffffff", -- 1e1a0
		x"ffffffff", -- 1e1a4
		x"ffffffff", -- 1e1a8
		x"ffffffff", -- 1e1ac
		x"ffffffff", -- 1e1b0
		x"ffffffff", -- 1e1b4
		x"ffffffff", -- 1e1b8
		x"ffffffff", -- 1e1bc
		x"ffffffff", -- 1e1c0
		x"ffffffff", -- 1e1c4
		x"ffffffff", -- 1e1c8
		x"ffffffff", -- 1e1cc
		x"ffffffff", -- 1e1d0
		x"ffffffff", -- 1e1d4
		x"ffffffff", -- 1e1d8
		x"ffffffff", -- 1e1dc
		x"ffffffff", -- 1e1e0
		x"ffffffff", -- 1e1e4
		x"ffffffff", -- 1e1e8
		x"ffffffff", -- 1e1ec
		x"ffffffff", -- 1e1f0
		x"ffffffff", -- 1e1f4
		x"ffffffff", -- 1e1f8
		x"ffffffff", -- 1e1fc
		x"ffffffff", -- 1e200
		x"ffffffff", -- 1e204
		x"ffffffff", -- 1e208
		x"ffffffff", -- 1e20c
		x"ffffffff", -- 1e210
		x"ffffffff", -- 1e214
		x"ffffffff", -- 1e218
		x"ffffffff", -- 1e21c
		x"ffffffff", -- 1e220
		x"ffffffff", -- 1e224
		x"ffffffff", -- 1e228
		x"ffffffff", -- 1e22c
		x"ffffffff", -- 1e230
		x"ffffffff", -- 1e234
		x"ffffffff", -- 1e238
		x"ffffffff", -- 1e23c
		x"ffffffff", -- 1e240
		x"ffffffff", -- 1e244
		x"ffffffff", -- 1e248
		x"ffffffff", -- 1e24c
		x"ffffffff", -- 1e250
		x"ffffffff", -- 1e254
		x"ffffffff", -- 1e258
		x"ffffffff", -- 1e25c
		x"ffffffff", -- 1e260
		x"ffffffff", -- 1e264
		x"ffffffff", -- 1e268
		x"ffffffff", -- 1e26c
		x"ffffffff", -- 1e270
		x"ffffffff", -- 1e274
		x"ffffffff", -- 1e278
		x"ffffffff", -- 1e27c
		x"ffffffff", -- 1e280
		x"ffffffff", -- 1e284
		x"ffffffff", -- 1e288
		x"ffffffff", -- 1e28c
		x"ffffffff", -- 1e290
		x"ffffffff", -- 1e294
		x"ffffffff", -- 1e298
		x"ffffffff", -- 1e29c
		x"ffffffff", -- 1e2a0
		x"ffffffff", -- 1e2a4
		x"ffffffff", -- 1e2a8
		x"ffffffff", -- 1e2ac
		x"ffffffff", -- 1e2b0
		x"ffffffff", -- 1e2b4
		x"ffffffff", -- 1e2b8
		x"ffffffff", -- 1e2bc
		x"ffffffff", -- 1e2c0
		x"ffffffff", -- 1e2c4
		x"ffffffff", -- 1e2c8
		x"ffffffff", -- 1e2cc
		x"ffffffff", -- 1e2d0
		x"ffffffff", -- 1e2d4
		x"ffffffff", -- 1e2d8
		x"ffffffff", -- 1e2dc
		x"ffffffff", -- 1e2e0
		x"ffffffff", -- 1e2e4
		x"ffffffff", -- 1e2e8
		x"ffffffff", -- 1e2ec
		x"ffffffff", -- 1e2f0
		x"ffffffff", -- 1e2f4
		x"ffffffff", -- 1e2f8
		x"ffffffff", -- 1e2fc
		x"ffffffff", -- 1e300
		x"ffffffff", -- 1e304
		x"ffffffff", -- 1e308
		x"ffffffff", -- 1e30c
		x"ffffffff", -- 1e310
		x"ffffffff", -- 1e314
		x"ffffffff", -- 1e318
		x"ffffffff", -- 1e31c
		x"ffffffff", -- 1e320
		x"ffffffff", -- 1e324
		x"ffffffff", -- 1e328
		x"ffffffff", -- 1e32c
		x"ffffffff", -- 1e330
		x"ffffffff", -- 1e334
		x"ffffffff", -- 1e338
		x"ffffffff", -- 1e33c
		x"ffffffff", -- 1e340
		x"ffffffff", -- 1e344
		x"ffffffff", -- 1e348
		x"ffffffff", -- 1e34c
		x"ffffffff", -- 1e350
		x"ffffffff", -- 1e354
		x"ffffffff", -- 1e358
		x"ffffffff", -- 1e35c
		x"ffffffff", -- 1e360
		x"ffffffff", -- 1e364
		x"ffffffff", -- 1e368
		x"ffffffff", -- 1e36c
		x"ffffffff", -- 1e370
		x"ffffffff", -- 1e374
		x"ffffffff", -- 1e378
		x"ffffffff", -- 1e37c
		x"ffffffff", -- 1e380
		x"ffffffff", -- 1e384
		x"ffffffff", -- 1e388
		x"ffffffff", -- 1e38c
		x"ffffffff", -- 1e390
		x"ffffffff", -- 1e394
		x"ffffffff", -- 1e398
		x"ffffffff", -- 1e39c
		x"ffffffff", -- 1e3a0
		x"ffffffff", -- 1e3a4
		x"ffffffff", -- 1e3a8
		x"ffffffff", -- 1e3ac
		x"ffffffff", -- 1e3b0
		x"ffffffff", -- 1e3b4
		x"ffffffff", -- 1e3b8
		x"ffffffff", -- 1e3bc
		x"ffffffff", -- 1e3c0
		x"ffffffff", -- 1e3c4
		x"ffffffff", -- 1e3c8
		x"ffffffff", -- 1e3cc
		x"ffffffff", -- 1e3d0
		x"ffffffff", -- 1e3d4
		x"ffffffff", -- 1e3d8
		x"ffffffff", -- 1e3dc
		x"ffffffff", -- 1e3e0
		x"ffffffff", -- 1e3e4
		x"ffffffff", -- 1e3e8
		x"ffffffff", -- 1e3ec
		x"ffffffff", -- 1e3f0
		x"ffffffff", -- 1e3f4
		x"ffffffff", -- 1e3f8
		x"ffffffff", -- 1e3fc
		x"ffffffff", -- 1e400
		x"ffffffff", -- 1e404
		x"ffffffff", -- 1e408
		x"ffffffff", -- 1e40c
		x"ffffffff", -- 1e410
		x"ffffffff", -- 1e414
		x"ffffffff", -- 1e418
		x"ffffffff", -- 1e41c
		x"ffffffff", -- 1e420
		x"ffffffff", -- 1e424
		x"ffffffff", -- 1e428
		x"ffffffff", -- 1e42c
		x"ffffffff", -- 1e430
		x"ffffffff", -- 1e434
		x"ffffffff", -- 1e438
		x"ffffffff", -- 1e43c
		x"ffffffff", -- 1e440
		x"ffffffff", -- 1e444
		x"ffffffff", -- 1e448
		x"ffffffff", -- 1e44c
		x"ffffffff", -- 1e450
		x"ffffffff", -- 1e454
		x"ffffffff", -- 1e458
		x"ffffffff", -- 1e45c
		x"ffffffff", -- 1e460
		x"ffffffff", -- 1e464
		x"ffffffff", -- 1e468
		x"ffffffff", -- 1e46c
		x"ffffffff", -- 1e470
		x"ffffffff", -- 1e474
		x"ffffffff", -- 1e478
		x"ffffffff", -- 1e47c
		x"ffffffff", -- 1e480
		x"ffffffff", -- 1e484
		x"ffffffff", -- 1e488
		x"ffffffff", -- 1e48c
		x"ffffffff", -- 1e490
		x"ffffffff", -- 1e494
		x"ffffffff", -- 1e498
		x"ffffffff", -- 1e49c
		x"ffffffff", -- 1e4a0
		x"ffffffff", -- 1e4a4
		x"ffffffff", -- 1e4a8
		x"ffffffff", -- 1e4ac
		x"ffffffff", -- 1e4b0
		x"ffffffff", -- 1e4b4
		x"ffffffff", -- 1e4b8
		x"ffffffff", -- 1e4bc
		x"ffffffff", -- 1e4c0
		x"ffffffff", -- 1e4c4
		x"ffffffff", -- 1e4c8
		x"ffffffff", -- 1e4cc
		x"ffffffff", -- 1e4d0
		x"ffffffff", -- 1e4d4
		x"ffffffff", -- 1e4d8
		x"ffffffff", -- 1e4dc
		x"ffffffff", -- 1e4e0
		x"ffffffff", -- 1e4e4
		x"ffffffff", -- 1e4e8
		x"ffffffff", -- 1e4ec
		x"ffffffff", -- 1e4f0
		x"ffffffff", -- 1e4f4
		x"ffffffff", -- 1e4f8
		x"ffffffff", -- 1e4fc
		x"ffffffff", -- 1e500
		x"ffffffff", -- 1e504
		x"ffffffff", -- 1e508
		x"ffffffff", -- 1e50c
		x"ffffffff", -- 1e510
		x"ffffffff", -- 1e514
		x"ffffffff", -- 1e518
		x"ffffffff", -- 1e51c
		x"ffffffff", -- 1e520
		x"ffffffff", -- 1e524
		x"ffffffff", -- 1e528
		x"ffffffff", -- 1e52c
		x"ffffffff", -- 1e530
		x"ffffffff", -- 1e534
		x"ffffffff", -- 1e538
		x"ffffffff", -- 1e53c
		x"ffffffff", -- 1e540
		x"ffffffff", -- 1e544
		x"ffffffff", -- 1e548
		x"ffffffff", -- 1e54c
		x"ffffffff", -- 1e550
		x"ffffffff", -- 1e554
		x"ffffffff", -- 1e558
		x"ffffffff", -- 1e55c
		x"ffffffff", -- 1e560
		x"ffffffff", -- 1e564
		x"ffffffff", -- 1e568
		x"ffffffff", -- 1e56c
		x"ffffffff", -- 1e570
		x"ffffffff", -- 1e574
		x"ffffffff", -- 1e578
		x"ffffffff", -- 1e57c
		x"ffffffff", -- 1e580
		x"ffffffff", -- 1e584
		x"ffffffff", -- 1e588
		x"ffffffff", -- 1e58c
		x"ffffffff", -- 1e590
		x"ffffffff", -- 1e594
		x"ffffffff", -- 1e598
		x"ffffffff", -- 1e59c
		x"ffffffff", -- 1e5a0
		x"ffffffff", -- 1e5a4
		x"ffffffff", -- 1e5a8
		x"ffffffff", -- 1e5ac
		x"ffffffff", -- 1e5b0
		x"ffffffff", -- 1e5b4
		x"ffffffff", -- 1e5b8
		x"ffffffff", -- 1e5bc
		x"ffffffff", -- 1e5c0
		x"ffffffff", -- 1e5c4
		x"ffffffff", -- 1e5c8
		x"ffffffff", -- 1e5cc
		x"ffffffff", -- 1e5d0
		x"ffffffff", -- 1e5d4
		x"ffffffff", -- 1e5d8
		x"ffffffff", -- 1e5dc
		x"ffffffff", -- 1e5e0
		x"ffffffff", -- 1e5e4
		x"ffffffff", -- 1e5e8
		x"ffffffff", -- 1e5ec
		x"ffffffff", -- 1e5f0
		x"ffffffff", -- 1e5f4
		x"ffffffff", -- 1e5f8
		x"ffffffff", -- 1e5fc
		x"ffffffff", -- 1e600
		x"ffffffff", -- 1e604
		x"ffffffff", -- 1e608
		x"ffffffff", -- 1e60c
		x"ffffffff", -- 1e610
		x"ffffffff", -- 1e614
		x"ffffffff", -- 1e618
		x"ffffffff", -- 1e61c
		x"ffffffff", -- 1e620
		x"ffffffff", -- 1e624
		x"ffffffff", -- 1e628
		x"ffffffff", -- 1e62c
		x"ffffffff", -- 1e630
		x"ffffffff", -- 1e634
		x"ffffffff", -- 1e638
		x"ffffffff", -- 1e63c
		x"ffffffff", -- 1e640
		x"ffffffff", -- 1e644
		x"ffffffff", -- 1e648
		x"ffffffff", -- 1e64c
		x"ffffffff", -- 1e650
		x"ffffffff", -- 1e654
		x"ffffffff", -- 1e658
		x"ffffffff", -- 1e65c
		x"ffffffff", -- 1e660
		x"ffffffff", -- 1e664
		x"ffffffff", -- 1e668
		x"ffffffff", -- 1e66c
		x"ffffffff", -- 1e670
		x"ffffffff", -- 1e674
		x"ffffffff", -- 1e678
		x"ffffffff", -- 1e67c
		x"ffffffff", -- 1e680
		x"ffffffff", -- 1e684
		x"ffffffff", -- 1e688
		x"ffffffff", -- 1e68c
		x"ffffffff", -- 1e690
		x"ffffffff", -- 1e694
		x"ffffffff", -- 1e698
		x"ffffffff", -- 1e69c
		x"ffffffff", -- 1e6a0
		x"ffffffff", -- 1e6a4
		x"ffffffff", -- 1e6a8
		x"ffffffff", -- 1e6ac
		x"ffffffff", -- 1e6b0
		x"ffffffff", -- 1e6b4
		x"ffffffff", -- 1e6b8
		x"ffffffff", -- 1e6bc
		x"ffffffff", -- 1e6c0
		x"ffffffff", -- 1e6c4
		x"ffffffff", -- 1e6c8
		x"ffffffff", -- 1e6cc
		x"ffffffff", -- 1e6d0
		x"ffffffff", -- 1e6d4
		x"ffffffff", -- 1e6d8
		x"ffffffff", -- 1e6dc
		x"ffffffff", -- 1e6e0
		x"ffffffff", -- 1e6e4
		x"ffffffff", -- 1e6e8
		x"ffffffff", -- 1e6ec
		x"ffffffff", -- 1e6f0
		x"ffffffff", -- 1e6f4
		x"ffffffff", -- 1e6f8
		x"ffffffff", -- 1e6fc
		x"ffffffff", -- 1e700
		x"ffffffff", -- 1e704
		x"ffffffff", -- 1e708
		x"ffffffff", -- 1e70c
		x"ffffffff", -- 1e710
		x"ffffffff", -- 1e714
		x"ffffffff", -- 1e718
		x"ffffffff", -- 1e71c
		x"ffffffff", -- 1e720
		x"ffffffff", -- 1e724
		x"ffffffff", -- 1e728
		x"ffffffff", -- 1e72c
		x"ffffffff", -- 1e730
		x"ffffffff", -- 1e734
		x"ffffffff", -- 1e738
		x"ffffffff", -- 1e73c
		x"ffffffff", -- 1e740
		x"ffffffff", -- 1e744
		x"ffffffff", -- 1e748
		x"ffffffff", -- 1e74c
		x"ffffffff", -- 1e750
		x"ffffffff", -- 1e754
		x"ffffffff", -- 1e758
		x"ffffffff", -- 1e75c
		x"ffffffff", -- 1e760
		x"ffffffff", -- 1e764
		x"ffffffff", -- 1e768
		x"ffffffff", -- 1e76c
		x"ffffffff", -- 1e770
		x"ffffffff", -- 1e774
		x"ffffffff", -- 1e778
		x"ffffffff", -- 1e77c
		x"ffffffff", -- 1e780
		x"ffffffff", -- 1e784
		x"ffffffff", -- 1e788
		x"ffffffff", -- 1e78c
		x"ffffffff", -- 1e790
		x"ffffffff", -- 1e794
		x"ffffffff", -- 1e798
		x"ffffffff", -- 1e79c
		x"ffffffff", -- 1e7a0
		x"ffffffff", -- 1e7a4
		x"ffffffff", -- 1e7a8
		x"ffffffff", -- 1e7ac
		x"ffffffff", -- 1e7b0
		x"ffffffff", -- 1e7b4
		x"ffffffff", -- 1e7b8
		x"ffffffff", -- 1e7bc
		x"ffffffff", -- 1e7c0
		x"ffffffff", -- 1e7c4
		x"ffffffff", -- 1e7c8
		x"ffffffff", -- 1e7cc
		x"ffffffff", -- 1e7d0
		x"ffffffff", -- 1e7d4
		x"ffffffff", -- 1e7d8
		x"ffffffff", -- 1e7dc
		x"ffffffff", -- 1e7e0
		x"ffffffff", -- 1e7e4
		x"ffffffff", -- 1e7e8
		x"ffffffff", -- 1e7ec
		x"ffffffff", -- 1e7f0
		x"ffffffff", -- 1e7f4
		x"ffffffff", -- 1e7f8
		x"ffffffff", -- 1e7fc
		x"ffffffff", -- 1e800
		x"ffffffff", -- 1e804
		x"ffffffff", -- 1e808
		x"ffffffff", -- 1e80c
		x"ffffffff", -- 1e810
		x"ffffffff", -- 1e814
		x"ffffffff", -- 1e818
		x"ffffffff", -- 1e81c
		x"ffffffff", -- 1e820
		x"ffffffff", -- 1e824
		x"ffffffff", -- 1e828
		x"ffffffff", -- 1e82c
		x"ffffffff", -- 1e830
		x"ffffffff", -- 1e834
		x"ffffffff", -- 1e838
		x"ffffffff", -- 1e83c
		x"ffffffff", -- 1e840
		x"ffffffff", -- 1e844
		x"ffffffff", -- 1e848
		x"ffffffff", -- 1e84c
		x"ffffffff", -- 1e850
		x"ffffffff", -- 1e854
		x"ffffffff", -- 1e858
		x"ffffffff", -- 1e85c
		x"ffffffff", -- 1e860
		x"ffffffff", -- 1e864
		x"ffffffff", -- 1e868
		x"ffffffff", -- 1e86c
		x"ffffffff", -- 1e870
		x"ffffffff", -- 1e874
		x"ffffffff", -- 1e878
		x"ffffffff", -- 1e87c
		x"ffffffff", -- 1e880
		x"ffffffff", -- 1e884
		x"ffffffff", -- 1e888
		x"ffffffff", -- 1e88c
		x"ffffffff", -- 1e890
		x"ffffffff", -- 1e894
		x"ffffffff", -- 1e898
		x"ffffffff", -- 1e89c
		x"ffffffff", -- 1e8a0
		x"ffffffff", -- 1e8a4
		x"ffffffff", -- 1e8a8
		x"ffffffff", -- 1e8ac
		x"ffffffff", -- 1e8b0
		x"ffffffff", -- 1e8b4
		x"ffffffff", -- 1e8b8
		x"ffffffff", -- 1e8bc
		x"ffffffff", -- 1e8c0
		x"ffffffff", -- 1e8c4
		x"ffffffff", -- 1e8c8
		x"ffffffff", -- 1e8cc
		x"ffffffff", -- 1e8d0
		x"ffffffff", -- 1e8d4
		x"ffffffff", -- 1e8d8
		x"ffffffff", -- 1e8dc
		x"ffffffff", -- 1e8e0
		x"ffffffff", -- 1e8e4
		x"ffffffff", -- 1e8e8
		x"ffffffff", -- 1e8ec
		x"ffffffff", -- 1e8f0
		x"ffffffff", -- 1e8f4
		x"ffffffff", -- 1e8f8
		x"ffffffff", -- 1e8fc
		x"ffffffff", -- 1e900
		x"ffffffff", -- 1e904
		x"ffffffff", -- 1e908
		x"ffffffff", -- 1e90c
		x"ffffffff", -- 1e910
		x"ffffffff", -- 1e914
		x"ffffffff", -- 1e918
		x"ffffffff", -- 1e91c
		x"ffffffff", -- 1e920
		x"ffffffff", -- 1e924
		x"ffffffff", -- 1e928
		x"ffffffff", -- 1e92c
		x"ffffffff", -- 1e930
		x"ffffffff", -- 1e934
		x"ffffffff", -- 1e938
		x"ffffffff", -- 1e93c
		x"ffffffff", -- 1e940
		x"ffffffff", -- 1e944
		x"ffffffff", -- 1e948
		x"ffffffff", -- 1e94c
		x"ffffffff", -- 1e950
		x"ffffffff", -- 1e954
		x"ffffffff", -- 1e958
		x"ffffffff", -- 1e95c
		x"ffffffff", -- 1e960
		x"ffffffff", -- 1e964
		x"ffffffff", -- 1e968
		x"ffffffff", -- 1e96c
		x"ffffffff", -- 1e970
		x"ffffffff", -- 1e974
		x"ffffffff", -- 1e978
		x"ffffffff", -- 1e97c
		x"ffffffff", -- 1e980
		x"ffffffff", -- 1e984
		x"ffffffff", -- 1e988
		x"ffffffff", -- 1e98c
		x"ffffffff", -- 1e990
		x"ffffffff", -- 1e994
		x"ffffffff", -- 1e998
		x"ffffffff", -- 1e99c
		x"ffffffff", -- 1e9a0
		x"ffffffff", -- 1e9a4
		x"ffffffff", -- 1e9a8
		x"ffffffff", -- 1e9ac
		x"ffffffff", -- 1e9b0
		x"ffffffff", -- 1e9b4
		x"ffffffff", -- 1e9b8
		x"ffffffff", -- 1e9bc
		x"ffffffff", -- 1e9c0
		x"ffffffff", -- 1e9c4
		x"ffffffff", -- 1e9c8
		x"ffffffff", -- 1e9cc
		x"ffffffff", -- 1e9d0
		x"ffffffff", -- 1e9d4
		x"ffffffff", -- 1e9d8
		x"ffffffff", -- 1e9dc
		x"ffffffff", -- 1e9e0
		x"ffffffff", -- 1e9e4
		x"ffffffff", -- 1e9e8
		x"ffffffff", -- 1e9ec
		x"ffffffff", -- 1e9f0
		x"ffffffff", -- 1e9f4
		x"ffffffff", -- 1e9f8
		x"ffffffff", -- 1e9fc
		x"ffffffff", -- 1ea00
		x"ffffffff", -- 1ea04
		x"ffffffff", -- 1ea08
		x"ffffffff", -- 1ea0c
		x"ffffffff", -- 1ea10
		x"ffffffff", -- 1ea14
		x"ffffffff", -- 1ea18
		x"ffffffff", -- 1ea1c
		x"ffffffff", -- 1ea20
		x"ffffffff", -- 1ea24
		x"ffffffff", -- 1ea28
		x"ffffffff", -- 1ea2c
		x"ffffffff", -- 1ea30
		x"ffffffff", -- 1ea34
		x"ffffffff", -- 1ea38
		x"ffffffff", -- 1ea3c
		x"ffffffff", -- 1ea40
		x"ffffffff", -- 1ea44
		x"ffffffff", -- 1ea48
		x"ffffffff", -- 1ea4c
		x"ffffffff", -- 1ea50
		x"ffffffff", -- 1ea54
		x"ffffffff", -- 1ea58
		x"ffffffff", -- 1ea5c
		x"ffffffff", -- 1ea60
		x"ffffffff", -- 1ea64
		x"ffffffff", -- 1ea68
		x"ffffffff", -- 1ea6c
		x"ffffffff", -- 1ea70
		x"ffffffff", -- 1ea74
		x"ffffffff", -- 1ea78
		x"ffffffff", -- 1ea7c
		x"ffffffff", -- 1ea80
		x"ffffffff", -- 1ea84
		x"ffffffff", -- 1ea88
		x"ffffffff", -- 1ea8c
		x"ffffffff", -- 1ea90
		x"ffffffff", -- 1ea94
		x"ffffffff", -- 1ea98
		x"ffffffff", -- 1ea9c
		x"ffffffff", -- 1eaa0
		x"ffffffff", -- 1eaa4
		x"ffffffff", -- 1eaa8
		x"ffffffff", -- 1eaac
		x"ffffffff", -- 1eab0
		x"ffffffff", -- 1eab4
		x"ffffffff", -- 1eab8
		x"ffffffff", -- 1eabc
		x"ffffffff", -- 1eac0
		x"ffffffff", -- 1eac4
		x"ffffffff", -- 1eac8
		x"ffffffff", -- 1eacc
		x"ffffffff", -- 1ead0
		x"ffffffff", -- 1ead4
		x"ffffffff", -- 1ead8
		x"ffffffff", -- 1eadc
		x"ffffffff", -- 1eae0
		x"ffffffff", -- 1eae4
		x"ffffffff", -- 1eae8
		x"ffffffff", -- 1eaec
		x"ffffffff", -- 1eaf0
		x"ffffffff", -- 1eaf4
		x"ffffffff", -- 1eaf8
		x"ffffffff", -- 1eafc
		x"ffffffff", -- 1eb00
		x"ffffffff", -- 1eb04
		x"ffffffff", -- 1eb08
		x"ffffffff", -- 1eb0c
		x"ffffffff", -- 1eb10
		x"ffffffff", -- 1eb14
		x"ffffffff", -- 1eb18
		x"ffffffff", -- 1eb1c
		x"ffffffff", -- 1eb20
		x"ffffffff", -- 1eb24
		x"ffffffff", -- 1eb28
		x"ffffffff", -- 1eb2c
		x"ffffffff", -- 1eb30
		x"ffffffff", -- 1eb34
		x"ffffffff", -- 1eb38
		x"ffffffff", -- 1eb3c
		x"ffffffff", -- 1eb40
		x"ffffffff", -- 1eb44
		x"ffffffff", -- 1eb48
		x"ffffffff", -- 1eb4c
		x"ffffffff", -- 1eb50
		x"ffffffff", -- 1eb54
		x"ffffffff", -- 1eb58
		x"ffffffff", -- 1eb5c
		x"ffffffff", -- 1eb60
		x"ffffffff", -- 1eb64
		x"ffffffff", -- 1eb68
		x"ffffffff", -- 1eb6c
		x"ffffffff", -- 1eb70
		x"ffffffff", -- 1eb74
		x"ffffffff", -- 1eb78
		x"ffffffff", -- 1eb7c
		x"ffffffff", -- 1eb80
		x"ffffffff", -- 1eb84
		x"ffffffff", -- 1eb88
		x"ffffffff", -- 1eb8c
		x"ffffffff", -- 1eb90
		x"ffffffff", -- 1eb94
		x"ffffffff", -- 1eb98
		x"ffffffff", -- 1eb9c
		x"ffffffff", -- 1eba0
		x"ffffffff", -- 1eba4
		x"ffffffff", -- 1eba8
		x"ffffffff", -- 1ebac
		x"ffffffff", -- 1ebb0
		x"ffffffff", -- 1ebb4
		x"ffffffff", -- 1ebb8
		x"ffffffff", -- 1ebbc
		x"ffffffff", -- 1ebc0
		x"ffffffff", -- 1ebc4
		x"ffffffff", -- 1ebc8
		x"ffffffff", -- 1ebcc
		x"ffffffff", -- 1ebd0
		x"ffffffff", -- 1ebd4
		x"ffffffff", -- 1ebd8
		x"ffffffff", -- 1ebdc
		x"ffffffff", -- 1ebe0
		x"ffffffff", -- 1ebe4
		x"ffffffff", -- 1ebe8
		x"ffffffff", -- 1ebec
		x"ffffffff", -- 1ebf0
		x"ffffffff", -- 1ebf4
		x"ffffffff", -- 1ebf8
		x"ffffffff", -- 1ebfc
		x"ffffffff", -- 1ec00
		x"ffffffff", -- 1ec04
		x"ffffffff", -- 1ec08
		x"ffffffff", -- 1ec0c
		x"ffffffff", -- 1ec10
		x"ffffffff", -- 1ec14
		x"ffffffff", -- 1ec18
		x"ffffffff", -- 1ec1c
		x"ffffffff", -- 1ec20
		x"ffffffff", -- 1ec24
		x"ffffffff", -- 1ec28
		x"ffffffff", -- 1ec2c
		x"ffffffff", -- 1ec30
		x"ffffffff", -- 1ec34
		x"ffffffff", -- 1ec38
		x"ffffffff", -- 1ec3c
		x"ffffffff", -- 1ec40
		x"ffffffff", -- 1ec44
		x"ffffffff", -- 1ec48
		x"ffffffff", -- 1ec4c
		x"ffffffff", -- 1ec50
		x"ffffffff", -- 1ec54
		x"ffffffff", -- 1ec58
		x"ffffffff", -- 1ec5c
		x"ffffffff", -- 1ec60
		x"ffffffff", -- 1ec64
		x"ffffffff", -- 1ec68
		x"ffffffff", -- 1ec6c
		x"ffffffff", -- 1ec70
		x"ffffffff", -- 1ec74
		x"ffffffff", -- 1ec78
		x"ffffffff", -- 1ec7c
		x"ffffffff", -- 1ec80
		x"ffffffff", -- 1ec84
		x"ffffffff", -- 1ec88
		x"ffffffff", -- 1ec8c
		x"ffffffff", -- 1ec90
		x"ffffffff", -- 1ec94
		x"ffffffff", -- 1ec98
		x"ffffffff", -- 1ec9c
		x"ffffffff", -- 1eca0
		x"ffffffff", -- 1eca4
		x"ffffffff", -- 1eca8
		x"ffffffff", -- 1ecac
		x"ffffffff", -- 1ecb0
		x"ffffffff", -- 1ecb4
		x"ffffffff", -- 1ecb8
		x"ffffffff", -- 1ecbc
		x"ffffffff", -- 1ecc0
		x"ffffffff", -- 1ecc4
		x"ffffffff", -- 1ecc8
		x"ffffffff", -- 1eccc
		x"ffffffff", -- 1ecd0
		x"ffffffff", -- 1ecd4
		x"ffffffff", -- 1ecd8
		x"ffffffff", -- 1ecdc
		x"ffffffff", -- 1ece0
		x"ffffffff", -- 1ece4
		x"ffffffff", -- 1ece8
		x"ffffffff", -- 1ecec
		x"ffffffff", -- 1ecf0
		x"ffffffff", -- 1ecf4
		x"ffffffff", -- 1ecf8
		x"ffffffff", -- 1ecfc
		x"ffffffff", -- 1ed00
		x"ffffffff", -- 1ed04
		x"ffffffff", -- 1ed08
		x"ffffffff", -- 1ed0c
		x"ffffffff", -- 1ed10
		x"ffffffff", -- 1ed14
		x"ffffffff", -- 1ed18
		x"ffffffff", -- 1ed1c
		x"ffffffff", -- 1ed20
		x"ffffffff", -- 1ed24
		x"ffffffff", -- 1ed28
		x"ffffffff", -- 1ed2c
		x"ffffffff", -- 1ed30
		x"ffffffff", -- 1ed34
		x"ffffffff", -- 1ed38
		x"ffffffff", -- 1ed3c
		x"ffffffff", -- 1ed40
		x"ffffffff", -- 1ed44
		x"ffffffff", -- 1ed48
		x"ffffffff", -- 1ed4c
		x"ffffffff", -- 1ed50
		x"ffffffff", -- 1ed54
		x"ffffffff", -- 1ed58
		x"ffffffff", -- 1ed5c
		x"ffffffff", -- 1ed60
		x"ffffffff", -- 1ed64
		x"ffffffff", -- 1ed68
		x"ffffffff", -- 1ed6c
		x"ffffffff", -- 1ed70
		x"ffffffff", -- 1ed74
		x"ffffffff", -- 1ed78
		x"ffffffff", -- 1ed7c
		x"ffffffff", -- 1ed80
		x"ffffffff", -- 1ed84
		x"ffffffff", -- 1ed88
		x"ffffffff", -- 1ed8c
		x"ffffffff", -- 1ed90
		x"ffffffff", -- 1ed94
		x"ffffffff", -- 1ed98
		x"ffffffff", -- 1ed9c
		x"ffffffff", -- 1eda0
		x"ffffffff", -- 1eda4
		x"ffffffff", -- 1eda8
		x"ffffffff", -- 1edac
		x"ffffffff", -- 1edb0
		x"ffffffff", -- 1edb4
		x"ffffffff", -- 1edb8
		x"ffffffff", -- 1edbc
		x"ffffffff", -- 1edc0
		x"ffffffff", -- 1edc4
		x"ffffffff", -- 1edc8
		x"ffffffff", -- 1edcc
		x"ffffffff", -- 1edd0
		x"ffffffff", -- 1edd4
		x"ffffffff", -- 1edd8
		x"ffffffff", -- 1eddc
		x"ffffffff", -- 1ede0
		x"ffffffff", -- 1ede4
		x"ffffffff", -- 1ede8
		x"ffffffff", -- 1edec
		x"ffffffff", -- 1edf0
		x"ffffffff", -- 1edf4
		x"ffffffff", -- 1edf8
		x"ffffffff", -- 1edfc
		x"ffffffff", -- 1ee00
		x"ffffffff", -- 1ee04
		x"ffffffff", -- 1ee08
		x"ffffffff", -- 1ee0c
		x"ffffffff", -- 1ee10
		x"ffffffff", -- 1ee14
		x"ffffffff", -- 1ee18
		x"ffffffff", -- 1ee1c
		x"ffffffff", -- 1ee20
		x"ffffffff", -- 1ee24
		x"ffffffff", -- 1ee28
		x"ffffffff", -- 1ee2c
		x"ffffffff", -- 1ee30
		x"ffffffff", -- 1ee34
		x"ffffffff", -- 1ee38
		x"ffffffff", -- 1ee3c
		x"ffffffff", -- 1ee40
		x"ffffffff", -- 1ee44
		x"ffffffff", -- 1ee48
		x"ffffffff", -- 1ee4c
		x"ffffffff", -- 1ee50
		x"ffffffff", -- 1ee54
		x"ffffffff", -- 1ee58
		x"ffffffff", -- 1ee5c
		x"ffffffff", -- 1ee60
		x"ffffffff", -- 1ee64
		x"ffffffff", -- 1ee68
		x"ffffffff", -- 1ee6c
		x"ffffffff", -- 1ee70
		x"ffffffff", -- 1ee74
		x"ffffffff", -- 1ee78
		x"ffffffff", -- 1ee7c
		x"ffffffff", -- 1ee80
		x"ffffffff", -- 1ee84
		x"ffffffff", -- 1ee88
		x"ffffffff", -- 1ee8c
		x"ffffffff", -- 1ee90
		x"ffffffff", -- 1ee94
		x"ffffffff", -- 1ee98
		x"ffffffff", -- 1ee9c
		x"ffffffff", -- 1eea0
		x"ffffffff", -- 1eea4
		x"ffffffff", -- 1eea8
		x"ffffffff", -- 1eeac
		x"ffffffff", -- 1eeb0
		x"ffffffff", -- 1eeb4
		x"ffffffff", -- 1eeb8
		x"ffffffff", -- 1eebc
		x"ffffffff", -- 1eec0
		x"ffffffff", -- 1eec4
		x"ffffffff", -- 1eec8
		x"ffffffff", -- 1eecc
		x"ffffffff", -- 1eed0
		x"ffffffff", -- 1eed4
		x"ffffffff", -- 1eed8
		x"ffffffff", -- 1eedc
		x"ffffffff", -- 1eee0
		x"ffffffff", -- 1eee4
		x"ffffffff", -- 1eee8
		x"ffffffff", -- 1eeec
		x"ffffffff", -- 1eef0
		x"ffffffff", -- 1eef4
		x"ffffffff", -- 1eef8
		x"ffffffff", -- 1eefc
		x"ffffffff", -- 1ef00
		x"ffffffff", -- 1ef04
		x"ffffffff", -- 1ef08
		x"ffffffff", -- 1ef0c
		x"ffffffff", -- 1ef10
		x"ffffffff", -- 1ef14
		x"ffffffff", -- 1ef18
		x"ffffffff", -- 1ef1c
		x"ffffffff", -- 1ef20
		x"ffffffff", -- 1ef24
		x"ffffffff", -- 1ef28
		x"ffffffff", -- 1ef2c
		x"ffffffff", -- 1ef30
		x"ffffffff", -- 1ef34
		x"ffffffff", -- 1ef38
		x"ffffffff", -- 1ef3c
		x"ffffffff", -- 1ef40
		x"ffffffff", -- 1ef44
		x"ffffffff", -- 1ef48
		x"ffffffff", -- 1ef4c
		x"ffffffff", -- 1ef50
		x"ffffffff", -- 1ef54
		x"ffffffff", -- 1ef58
		x"ffffffff", -- 1ef5c
		x"ffffffff", -- 1ef60
		x"ffffffff", -- 1ef64
		x"ffffffff", -- 1ef68
		x"ffffffff", -- 1ef6c
		x"ffffffff", -- 1ef70
		x"ffffffff", -- 1ef74
		x"ffffffff", -- 1ef78
		x"ffffffff", -- 1ef7c
		x"ffffffff", -- 1ef80
		x"ffffffff", -- 1ef84
		x"ffffffff", -- 1ef88
		x"ffffffff", -- 1ef8c
		x"ffffffff", -- 1ef90
		x"ffffffff", -- 1ef94
		x"ffffffff", -- 1ef98
		x"ffffffff", -- 1ef9c
		x"ffffffff", -- 1efa0
		x"ffffffff", -- 1efa4
		x"ffffffff", -- 1efa8
		x"ffffffff", -- 1efac
		x"ffffffff", -- 1efb0
		x"ffffffff", -- 1efb4
		x"ffffffff", -- 1efb8
		x"ffffffff", -- 1efbc
		x"ffffffff", -- 1efc0
		x"ffffffff", -- 1efc4
		x"ffffffff", -- 1efc8
		x"ffffffff", -- 1efcc
		x"ffffffff", -- 1efd0
		x"ffffffff", -- 1efd4
		x"ffffffff", -- 1efd8
		x"ffffffff", -- 1efdc
		x"ffffffff", -- 1efe0
		x"ffffffff", -- 1efe4
		x"ffffffff", -- 1efe8
		x"ffffffff", -- 1efec
		x"ffffffff", -- 1eff0
		x"ffffffff", -- 1eff4
		x"ffffffff", -- 1eff8
		x"ffffffff", -- 1effc
		x"ffffffff", -- 1f000
		x"ffffffff", -- 1f004
		x"ffffffff", -- 1f008
		x"ffffffff", -- 1f00c
		x"ffffffff", -- 1f010
		x"ffffffff", -- 1f014
		x"ffffffff", -- 1f018
		x"ffffffff", -- 1f01c
		x"ffffffff", -- 1f020
		x"ffffffff", -- 1f024
		x"ffffffff", -- 1f028
		x"ffffffff", -- 1f02c
		x"ffffffff", -- 1f030
		x"ffffffff", -- 1f034
		x"ffffffff", -- 1f038
		x"ffffffff", -- 1f03c
		x"ffffffff", -- 1f040
		x"ffffffff", -- 1f044
		x"ffffffff", -- 1f048
		x"ffffffff", -- 1f04c
		x"ffffffff", -- 1f050
		x"ffffffff", -- 1f054
		x"ffffffff", -- 1f058
		x"ffffffff", -- 1f05c
		x"ffffffff", -- 1f060
		x"ffffffff", -- 1f064
		x"ffffffff", -- 1f068
		x"ffffffff", -- 1f06c
		x"ffffffff", -- 1f070
		x"ffffffff", -- 1f074
		x"ffffffff", -- 1f078
		x"ffffffff", -- 1f07c
		x"ffffffff", -- 1f080
		x"ffffffff", -- 1f084
		x"ffffffff", -- 1f088
		x"ffffffff", -- 1f08c
		x"ffffffff", -- 1f090
		x"ffffffff", -- 1f094
		x"ffffffff", -- 1f098
		x"ffffffff", -- 1f09c
		x"ffffffff", -- 1f0a0
		x"ffffffff", -- 1f0a4
		x"ffffffff", -- 1f0a8
		x"ffffffff", -- 1f0ac
		x"ffffffff", -- 1f0b0
		x"ffffffff", -- 1f0b4
		x"ffffffff", -- 1f0b8
		x"ffffffff", -- 1f0bc
		x"ffffffff", -- 1f0c0
		x"ffffffff", -- 1f0c4
		x"ffffffff", -- 1f0c8
		x"ffffffff", -- 1f0cc
		x"ffffffff", -- 1f0d0
		x"ffffffff", -- 1f0d4
		x"ffffffff", -- 1f0d8
		x"ffffffff", -- 1f0dc
		x"ffffffff", -- 1f0e0
		x"ffffffff", -- 1f0e4
		x"ffffffff", -- 1f0e8
		x"ffffffff", -- 1f0ec
		x"ffffffff", -- 1f0f0
		x"ffffffff", -- 1f0f4
		x"ffffffff", -- 1f0f8
		x"ffffffff", -- 1f0fc
		x"ffffffff", -- 1f100
		x"ffffffff", -- 1f104
		x"ffffffff", -- 1f108
		x"ffffffff", -- 1f10c
		x"ffffffff", -- 1f110
		x"ffffffff", -- 1f114
		x"ffffffff", -- 1f118
		x"ffffffff", -- 1f11c
		x"ffffffff", -- 1f120
		x"ffffffff", -- 1f124
		x"ffffffff", -- 1f128
		x"ffffffff", -- 1f12c
		x"ffffffff", -- 1f130
		x"ffffffff", -- 1f134
		x"ffffffff", -- 1f138
		x"ffffffff", -- 1f13c
		x"ffffffff", -- 1f140
		x"ffffffff", -- 1f144
		x"ffffffff", -- 1f148
		x"ffffffff", -- 1f14c
		x"ffffffff", -- 1f150
		x"ffffffff", -- 1f154
		x"ffffffff", -- 1f158
		x"ffffffff", -- 1f15c
		x"ffffffff", -- 1f160
		x"ffffffff", -- 1f164
		x"ffffffff", -- 1f168
		x"ffffffff", -- 1f16c
		x"ffffffff", -- 1f170
		x"ffffffff", -- 1f174
		x"ffffffff", -- 1f178
		x"ffffffff", -- 1f17c
		x"ffffffff", -- 1f180
		x"ffffffff", -- 1f184
		x"ffffffff", -- 1f188
		x"ffffffff", -- 1f18c
		x"ffffffff", -- 1f190
		x"ffffffff", -- 1f194
		x"ffffffff", -- 1f198
		x"ffffffff", -- 1f19c
		x"ffffffff", -- 1f1a0
		x"ffffffff", -- 1f1a4
		x"ffffffff", -- 1f1a8
		x"ffffffff", -- 1f1ac
		x"ffffffff", -- 1f1b0
		x"ffffffff", -- 1f1b4
		x"ffffffff", -- 1f1b8
		x"ffffffff", -- 1f1bc
		x"ffffffff", -- 1f1c0
		x"ffffffff", -- 1f1c4
		x"ffffffff", -- 1f1c8
		x"ffffffff", -- 1f1cc
		x"ffffffff", -- 1f1d0
		x"ffffffff", -- 1f1d4
		x"ffffffff", -- 1f1d8
		x"ffffffff", -- 1f1dc
		x"ffffffff", -- 1f1e0
		x"ffffffff", -- 1f1e4
		x"ffffffff", -- 1f1e8
		x"ffffffff", -- 1f1ec
		x"ffffffff", -- 1f1f0
		x"ffffffff", -- 1f1f4
		x"ffffffff", -- 1f1f8
		x"ffffffff", -- 1f1fc
		x"ffffffff", -- 1f200
		x"ffffffff", -- 1f204
		x"ffffffff", -- 1f208
		x"ffffffff", -- 1f20c
		x"ffffffff", -- 1f210
		x"ffffffff", -- 1f214
		x"ffffffff", -- 1f218
		x"ffffffff", -- 1f21c
		x"ffffffff", -- 1f220
		x"ffffffff", -- 1f224
		x"ffffffff", -- 1f228
		x"ffffffff", -- 1f22c
		x"ffffffff", -- 1f230
		x"ffffffff", -- 1f234
		x"ffffffff", -- 1f238
		x"ffffffff", -- 1f23c
		x"ffffffff", -- 1f240
		x"ffffffff", -- 1f244
		x"ffffffff", -- 1f248
		x"ffffffff", -- 1f24c
		x"ffffffff", -- 1f250
		x"ffffffff", -- 1f254
		x"ffffffff", -- 1f258
		x"ffffffff", -- 1f25c
		x"ffffffff", -- 1f260
		x"ffffffff", -- 1f264
		x"ffffffff", -- 1f268
		x"ffffffff", -- 1f26c
		x"ffffffff", -- 1f270
		x"ffffffff", -- 1f274
		x"ffffffff", -- 1f278
		x"ffffffff", -- 1f27c
		x"ffffffff", -- 1f280
		x"ffffffff", -- 1f284
		x"ffffffff", -- 1f288
		x"ffffffff", -- 1f28c
		x"ffffffff", -- 1f290
		x"ffffffff", -- 1f294
		x"ffffffff", -- 1f298
		x"ffffffff", -- 1f29c
		x"ffffffff", -- 1f2a0
		x"ffffffff", -- 1f2a4
		x"ffffffff", -- 1f2a8
		x"ffffffff", -- 1f2ac
		x"ffffffff", -- 1f2b0
		x"ffffffff", -- 1f2b4
		x"ffffffff", -- 1f2b8
		x"ffffffff", -- 1f2bc
		x"ffffffff", -- 1f2c0
		x"ffffffff", -- 1f2c4
		x"ffffffff", -- 1f2c8
		x"ffffffff", -- 1f2cc
		x"ffffffff", -- 1f2d0
		x"ffffffff", -- 1f2d4
		x"ffffffff", -- 1f2d8
		x"ffffffff", -- 1f2dc
		x"ffffffff", -- 1f2e0
		x"ffffffff", -- 1f2e4
		x"ffffffff", -- 1f2e8
		x"ffffffff", -- 1f2ec
		x"ffffffff", -- 1f2f0
		x"ffffffff", -- 1f2f4
		x"ffffffff", -- 1f2f8
		x"ffffffff", -- 1f2fc
		x"ffffffff", -- 1f300
		x"ffffffff", -- 1f304
		x"ffffffff", -- 1f308
		x"ffffffff", -- 1f30c
		x"ffffffff", -- 1f310
		x"ffffffff", -- 1f314
		x"ffffffff", -- 1f318
		x"ffffffff", -- 1f31c
		x"ffffffff", -- 1f320
		x"ffffffff", -- 1f324
		x"ffffffff", -- 1f328
		x"ffffffff", -- 1f32c
		x"ffffffff", -- 1f330
		x"ffffffff", -- 1f334
		x"ffffffff", -- 1f338
		x"ffffffff", -- 1f33c
		x"ffffffff", -- 1f340
		x"ffffffff", -- 1f344
		x"ffffffff", -- 1f348
		x"ffffffff", -- 1f34c
		x"ffffffff", -- 1f350
		x"ffffffff", -- 1f354
		x"ffffffff", -- 1f358
		x"ffffffff", -- 1f35c
		x"ffffffff", -- 1f360
		x"ffffffff", -- 1f364
		x"ffffffff", -- 1f368
		x"ffffffff", -- 1f36c
		x"ffffffff", -- 1f370
		x"ffffffff", -- 1f374
		x"ffffffff", -- 1f378
		x"ffffffff", -- 1f37c
		x"ffffffff", -- 1f380
		x"ffffffff", -- 1f384
		x"ffffffff", -- 1f388
		x"ffffffff", -- 1f38c
		x"ffffffff", -- 1f390
		x"ffffffff", -- 1f394
		x"ffffffff", -- 1f398
		x"ffffffff", -- 1f39c
		x"ffffffff", -- 1f3a0
		x"ffffffff", -- 1f3a4
		x"ffffffff", -- 1f3a8
		x"ffffffff", -- 1f3ac
		x"ffffffff", -- 1f3b0
		x"ffffffff", -- 1f3b4
		x"ffffffff", -- 1f3b8
		x"ffffffff", -- 1f3bc
		x"ffffffff", -- 1f3c0
		x"ffffffff", -- 1f3c4
		x"ffffffff", -- 1f3c8
		x"ffffffff", -- 1f3cc
		x"ffffffff", -- 1f3d0
		x"ffffffff", -- 1f3d4
		x"ffffffff", -- 1f3d8
		x"ffffffff", -- 1f3dc
		x"ffffffff", -- 1f3e0
		x"ffffffff", -- 1f3e4
		x"ffffffff", -- 1f3e8
		x"ffffffff", -- 1f3ec
		x"ffffffff", -- 1f3f0
		x"ffffffff", -- 1f3f4
		x"ffffffff", -- 1f3f8
		x"ffffffff", -- 1f3fc
		x"ffffffff", -- 1f400
		x"ffffffff", -- 1f404
		x"ffffffff", -- 1f408
		x"ffffffff", -- 1f40c
		x"ffffffff", -- 1f410
		x"ffffffff", -- 1f414
		x"ffffffff", -- 1f418
		x"ffffffff", -- 1f41c
		x"ffffffff", -- 1f420
		x"ffffffff", -- 1f424
		x"ffffffff", -- 1f428
		x"ffffffff", -- 1f42c
		x"ffffffff", -- 1f430
		x"ffffffff", -- 1f434
		x"ffffffff", -- 1f438
		x"ffffffff", -- 1f43c
		x"ffffffff", -- 1f440
		x"ffffffff", -- 1f444
		x"ffffffff", -- 1f448
		x"ffffffff", -- 1f44c
		x"ffffffff", -- 1f450
		x"ffffffff", -- 1f454
		x"ffffffff", -- 1f458
		x"ffffffff", -- 1f45c
		x"ffffffff", -- 1f460
		x"ffffffff", -- 1f464
		x"ffffffff", -- 1f468
		x"ffffffff", -- 1f46c
		x"ffffffff", -- 1f470
		x"ffffffff", -- 1f474
		x"ffffffff", -- 1f478
		x"ffffffff", -- 1f47c
		x"ffffffff", -- 1f480
		x"ffffffff", -- 1f484
		x"ffffffff", -- 1f488
		x"ffffffff", -- 1f48c
		x"ffffffff", -- 1f490
		x"ffffffff", -- 1f494
		x"ffffffff", -- 1f498
		x"ffffffff", -- 1f49c
		x"ffffffff", -- 1f4a0
		x"ffffffff", -- 1f4a4
		x"ffffffff", -- 1f4a8
		x"ffffffff", -- 1f4ac
		x"ffffffff", -- 1f4b0
		x"ffffffff", -- 1f4b4
		x"ffffffff", -- 1f4b8
		x"ffffffff", -- 1f4bc
		x"ffffffff", -- 1f4c0
		x"ffffffff", -- 1f4c4
		x"ffffffff", -- 1f4c8
		x"ffffffff", -- 1f4cc
		x"ffffffff", -- 1f4d0
		x"ffffffff", -- 1f4d4
		x"ffffffff", -- 1f4d8
		x"ffffffff", -- 1f4dc
		x"ffffffff", -- 1f4e0
		x"ffffffff", -- 1f4e4
		x"ffffffff", -- 1f4e8
		x"ffffffff", -- 1f4ec
		x"ffffffff", -- 1f4f0
		x"ffffffff", -- 1f4f4
		x"ffffffff", -- 1f4f8
		x"ffffffff", -- 1f4fc
		x"ffffffff", -- 1f500
		x"ffffffff", -- 1f504
		x"ffffffff", -- 1f508
		x"ffffffff", -- 1f50c
		x"ffffffff", -- 1f510
		x"ffffffff", -- 1f514
		x"ffffffff", -- 1f518
		x"ffffffff", -- 1f51c
		x"ffffffff", -- 1f520
		x"ffffffff", -- 1f524
		x"ffffffff", -- 1f528
		x"ffffffff", -- 1f52c
		x"ffffffff", -- 1f530
		x"ffffffff", -- 1f534
		x"ffffffff", -- 1f538
		x"ffffffff", -- 1f53c
		x"ffffffff", -- 1f540
		x"ffffffff", -- 1f544
		x"ffffffff", -- 1f548
		x"ffffffff", -- 1f54c
		x"ffffffff", -- 1f550
		x"ffffffff", -- 1f554
		x"ffffffff", -- 1f558
		x"ffffffff", -- 1f55c
		x"ffffffff", -- 1f560
		x"ffffffff", -- 1f564
		x"ffffffff", -- 1f568
		x"ffffffff", -- 1f56c
		x"ffffffff", -- 1f570
		x"ffffffff", -- 1f574
		x"ffffffff", -- 1f578
		x"ffffffff", -- 1f57c
		x"ffffffff", -- 1f580
		x"ffffffff", -- 1f584
		x"ffffffff", -- 1f588
		x"ffffffff", -- 1f58c
		x"ffffffff", -- 1f590
		x"ffffffff", -- 1f594
		x"ffffffff", -- 1f598
		x"ffffffff", -- 1f59c
		x"ffffffff", -- 1f5a0
		x"ffffffff", -- 1f5a4
		x"ffffffff", -- 1f5a8
		x"ffffffff", -- 1f5ac
		x"ffffffff", -- 1f5b0
		x"ffffffff", -- 1f5b4
		x"ffffffff", -- 1f5b8
		x"ffffffff", -- 1f5bc
		x"ffffffff", -- 1f5c0
		x"ffffffff", -- 1f5c4
		x"ffffffff", -- 1f5c8
		x"ffffffff", -- 1f5cc
		x"ffffffff", -- 1f5d0
		x"ffffffff", -- 1f5d4
		x"ffffffff", -- 1f5d8
		x"ffffffff", -- 1f5dc
		x"ffffffff", -- 1f5e0
		x"ffffffff", -- 1f5e4
		x"ffffffff", -- 1f5e8
		x"ffffffff", -- 1f5ec
		x"ffffffff", -- 1f5f0
		x"ffffffff", -- 1f5f4
		x"ffffffff", -- 1f5f8
		x"ffffffff", -- 1f5fc
		x"ffffffff", -- 1f600
		x"ffffffff", -- 1f604
		x"ffffffff", -- 1f608
		x"ffffffff", -- 1f60c
		x"ffffffff", -- 1f610
		x"ffffffff", -- 1f614
		x"ffffffff", -- 1f618
		x"ffffffff", -- 1f61c
		x"ffffffff", -- 1f620
		x"ffffffff", -- 1f624
		x"ffffffff", -- 1f628
		x"ffffffff", -- 1f62c
		x"ffffffff", -- 1f630
		x"ffffffff", -- 1f634
		x"ffffffff", -- 1f638
		x"ffffffff", -- 1f63c
		x"ffffffff", -- 1f640
		x"ffffffff", -- 1f644
		x"ffffffff", -- 1f648
		x"ffffffff", -- 1f64c
		x"ffffffff", -- 1f650
		x"ffffffff", -- 1f654
		x"ffffffff", -- 1f658
		x"ffffffff", -- 1f65c
		x"ffffffff", -- 1f660
		x"ffffffff", -- 1f664
		x"ffffffff", -- 1f668
		x"ffffffff", -- 1f66c
		x"ffffffff", -- 1f670
		x"ffffffff", -- 1f674
		x"ffffffff", -- 1f678
		x"ffffffff", -- 1f67c
		x"ffffffff", -- 1f680
		x"ffffffff", -- 1f684
		x"ffffffff", -- 1f688
		x"ffffffff", -- 1f68c
		x"ffffffff", -- 1f690
		x"ffffffff", -- 1f694
		x"ffffffff", -- 1f698
		x"ffffffff", -- 1f69c
		x"ffffffff", -- 1f6a0
		x"ffffffff", -- 1f6a4
		x"ffffffff", -- 1f6a8
		x"ffffffff", -- 1f6ac
		x"ffffffff", -- 1f6b0
		x"ffffffff", -- 1f6b4
		x"ffffffff", -- 1f6b8
		x"ffffffff", -- 1f6bc
		x"ffffffff", -- 1f6c0
		x"ffffffff", -- 1f6c4
		x"ffffffff", -- 1f6c8
		x"ffffffff", -- 1f6cc
		x"ffffffff", -- 1f6d0
		x"ffffffff", -- 1f6d4
		x"ffffffff", -- 1f6d8
		x"ffffffff", -- 1f6dc
		x"ffffffff", -- 1f6e0
		x"ffffffff", -- 1f6e4
		x"ffffffff", -- 1f6e8
		x"ffffffff", -- 1f6ec
		x"ffffffff", -- 1f6f0
		x"ffffffff", -- 1f6f4
		x"ffffffff", -- 1f6f8
		x"ffffffff", -- 1f6fc
		x"ffffffff", -- 1f700
		x"ffffffff", -- 1f704
		x"ffffffff", -- 1f708
		x"ffffffff", -- 1f70c
		x"ffffffff", -- 1f710
		x"ffffffff", -- 1f714
		x"ffffffff", -- 1f718
		x"ffffffff", -- 1f71c
		x"ffffffff", -- 1f720
		x"ffffffff", -- 1f724
		x"ffffffff", -- 1f728
		x"ffffffff", -- 1f72c
		x"ffffffff", -- 1f730
		x"ffffffff", -- 1f734
		x"ffffffff", -- 1f738
		x"ffffffff", -- 1f73c
		x"ffffffff", -- 1f740
		x"ffffffff", -- 1f744
		x"ffffffff", -- 1f748
		x"ffffffff", -- 1f74c
		x"ffffffff", -- 1f750
		x"ffffffff", -- 1f754
		x"ffffffff", -- 1f758
		x"ffffffff", -- 1f75c
		x"ffffffff", -- 1f760
		x"ffffffff", -- 1f764
		x"ffffffff", -- 1f768
		x"ffffffff", -- 1f76c
		x"ffffffff", -- 1f770
		x"ffffffff", -- 1f774
		x"ffffffff", -- 1f778
		x"ffffffff", -- 1f77c
		x"ffffffff", -- 1f780
		x"ffffffff", -- 1f784
		x"ffffffff", -- 1f788
		x"ffffffff", -- 1f78c
		x"ffffffff", -- 1f790
		x"ffffffff", -- 1f794
		x"ffffffff", -- 1f798
		x"ffffffff", -- 1f79c
		x"ffffffff", -- 1f7a0
		x"ffffffff", -- 1f7a4
		x"ffffffff", -- 1f7a8
		x"ffffffff", -- 1f7ac
		x"ffffffff", -- 1f7b0
		x"ffffffff", -- 1f7b4
		x"ffffffff", -- 1f7b8
		x"ffffffff", -- 1f7bc
		x"ffffffff", -- 1f7c0
		x"ffffffff", -- 1f7c4
		x"ffffffff", -- 1f7c8
		x"ffffffff", -- 1f7cc
		x"ffffffff", -- 1f7d0
		x"ffffffff", -- 1f7d4
		x"ffffffff", -- 1f7d8
		x"ffffffff", -- 1f7dc
		x"ffffffff", -- 1f7e0
		x"ffffffff", -- 1f7e4
		x"ffffffff", -- 1f7e8
		x"ffffffff", -- 1f7ec
		x"ffffffff", -- 1f7f0
		x"ffffffff", -- 1f7f4
		x"ffffffff", -- 1f7f8
		x"ffffffff", -- 1f7fc
		x"ffffffff", -- 1f800
		x"ffffffff", -- 1f804
		x"ffffffff", -- 1f808
		x"ffffffff", -- 1f80c
		x"ffffffff", -- 1f810
		x"ffffffff", -- 1f814
		x"ffffffff", -- 1f818
		x"ffffffff", -- 1f81c
		x"ffffffff", -- 1f820
		x"ffffffff", -- 1f824
		x"ffffffff", -- 1f828
		x"ffffffff", -- 1f82c
		x"ffffffff", -- 1f830
		x"ffffffff", -- 1f834
		x"ffffffff", -- 1f838
		x"ffffffff", -- 1f83c
		x"ffffffff", -- 1f840
		x"ffffffff", -- 1f844
		x"ffffffff", -- 1f848
		x"ffffffff", -- 1f84c
		x"ffffffff", -- 1f850
		x"ffffffff", -- 1f854
		x"ffffffff", -- 1f858
		x"ffffffff", -- 1f85c
		x"ffffffff", -- 1f860
		x"ffffffff", -- 1f864
		x"ffffffff", -- 1f868
		x"ffffffff", -- 1f86c
		x"ffffffff", -- 1f870
		x"ffffffff", -- 1f874
		x"ffffffff", -- 1f878
		x"ffffffff", -- 1f87c
		x"ffffffff", -- 1f880
		x"ffffffff", -- 1f884
		x"ffffffff", -- 1f888
		x"ffffffff", -- 1f88c
		x"ffffffff", -- 1f890
		x"ffffffff", -- 1f894
		x"ffffffff", -- 1f898
		x"ffffffff", -- 1f89c
		x"ffffffff", -- 1f8a0
		x"ffffffff", -- 1f8a4
		x"ffffffff", -- 1f8a8
		x"ffffffff", -- 1f8ac
		x"ffffffff", -- 1f8b0
		x"ffffffff", -- 1f8b4
		x"ffffffff", -- 1f8b8
		x"ffffffff", -- 1f8bc
		x"ffffffff", -- 1f8c0
		x"ffffffff", -- 1f8c4
		x"ffffffff", -- 1f8c8
		x"ffffffff", -- 1f8cc
		x"ffffffff", -- 1f8d0
		x"ffffffff", -- 1f8d4
		x"ffffffff", -- 1f8d8
		x"ffffffff", -- 1f8dc
		x"ffffffff", -- 1f8e0
		x"ffffffff", -- 1f8e4
		x"ffffffff", -- 1f8e8
		x"ffffffff", -- 1f8ec
		x"ffffffff", -- 1f8f0
		x"ffffffff", -- 1f8f4
		x"ffffffff", -- 1f8f8
		x"ffffffff", -- 1f8fc
		x"ffffffff", -- 1f900
		x"ffffffff", -- 1f904
		x"ffffffff", -- 1f908
		x"ffffffff", -- 1f90c
		x"ffffffff", -- 1f910
		x"ffffffff", -- 1f914
		x"ffffffff", -- 1f918
		x"ffffffff", -- 1f91c
		x"ffffffff", -- 1f920
		x"ffffffff", -- 1f924
		x"ffffffff", -- 1f928
		x"ffffffff", -- 1f92c
		x"ffffffff", -- 1f930
		x"ffffffff", -- 1f934
		x"ffffffff", -- 1f938
		x"ffffffff", -- 1f93c
		x"ffffffff", -- 1f940
		x"ffffffff", -- 1f944
		x"ffffffff", -- 1f948
		x"ffffffff", -- 1f94c
		x"ffffffff", -- 1f950
		x"ffffffff", -- 1f954
		x"ffffffff", -- 1f958
		x"ffffffff", -- 1f95c
		x"ffffffff", -- 1f960
		x"ffffffff", -- 1f964
		x"ffffffff", -- 1f968
		x"ffffffff", -- 1f96c
		x"ffffffff", -- 1f970
		x"ffffffff", -- 1f974
		x"ffffffff", -- 1f978
		x"ffffffff", -- 1f97c
		x"ffffffff", -- 1f980
		x"ffffffff", -- 1f984
		x"ffffffff", -- 1f988
		x"ffffffff", -- 1f98c
		x"ffffffff", -- 1f990
		x"ffffffff", -- 1f994
		x"ffffffff", -- 1f998
		x"ffffffff", -- 1f99c
		x"ffffffff", -- 1f9a0
		x"ffffffff", -- 1f9a4
		x"ffffffff", -- 1f9a8
		x"ffffffff", -- 1f9ac
		x"ffffffff", -- 1f9b0
		x"ffffffff", -- 1f9b4
		x"ffffffff", -- 1f9b8
		x"ffffffff", -- 1f9bc
		x"ffffffff", -- 1f9c0
		x"ffffffff", -- 1f9c4
		x"ffffffff", -- 1f9c8
		x"ffffffff", -- 1f9cc
		x"ffffffff", -- 1f9d0
		x"ffffffff", -- 1f9d4
		x"ffffffff", -- 1f9d8
		x"ffffffff", -- 1f9dc
		x"ffffffff", -- 1f9e0
		x"ffffffff", -- 1f9e4
		x"ffffffff", -- 1f9e8
		x"ffffffff", -- 1f9ec
		x"ffffffff", -- 1f9f0
		x"ffffffff", -- 1f9f4
		x"ffffffff", -- 1f9f8
		x"ffffffff", -- 1f9fc
		x"ffffffff", -- 1fa00
		x"ffffffff", -- 1fa04
		x"ffffffff", -- 1fa08
		x"ffffffff", -- 1fa0c
		x"ffffffff", -- 1fa10
		x"ffffffff", -- 1fa14
		x"ffffffff", -- 1fa18
		x"ffffffff", -- 1fa1c
		x"ffffffff", -- 1fa20
		x"ffffffff", -- 1fa24
		x"ffffffff", -- 1fa28
		x"ffffffff", -- 1fa2c
		x"ffffffff", -- 1fa30
		x"ffffffff", -- 1fa34
		x"ffffffff", -- 1fa38
		x"ffffffff", -- 1fa3c
		x"ffffffff", -- 1fa40
		x"ffffffff", -- 1fa44
		x"ffffffff", -- 1fa48
		x"ffffffff", -- 1fa4c
		x"ffffffff", -- 1fa50
		x"ffffffff", -- 1fa54
		x"ffffffff", -- 1fa58
		x"ffffffff", -- 1fa5c
		x"ffffffff", -- 1fa60
		x"ffffffff", -- 1fa64
		x"ffffffff", -- 1fa68
		x"ffffffff", -- 1fa6c
		x"ffffffff", -- 1fa70
		x"ffffffff", -- 1fa74
		x"ffffffff", -- 1fa78
		x"ffffffff", -- 1fa7c
		x"ffffffff", -- 1fa80
		x"ffffffff", -- 1fa84
		x"ffffffff", -- 1fa88
		x"ffffffff", -- 1fa8c
		x"ffffffff", -- 1fa90
		x"ffffffff", -- 1fa94
		x"ffffffff", -- 1fa98
		x"ffffffff", -- 1fa9c
		x"ffffffff", -- 1faa0
		x"ffffffff", -- 1faa4
		x"ffffffff", -- 1faa8
		x"ffffffff", -- 1faac
		x"ffffffff", -- 1fab0
		x"ffffffff", -- 1fab4
		x"ffffffff", -- 1fab8
		x"ffffffff", -- 1fabc
		x"ffffffff", -- 1fac0
		x"ffffffff", -- 1fac4
		x"ffffffff", -- 1fac8
		x"ffffffff", -- 1facc
		x"ffffffff", -- 1fad0
		x"ffffffff", -- 1fad4
		x"ffffffff", -- 1fad8
		x"ffffffff", -- 1fadc
		x"ffffffff", -- 1fae0
		x"ffffffff", -- 1fae4
		x"ffffffff", -- 1fae8
		x"ffffffff", -- 1faec
		x"ffffffff", -- 1faf0
		x"ffffffff", -- 1faf4
		x"ffffffff", -- 1faf8
		x"ffffffff", -- 1fafc
		x"ffffffff", -- 1fb00
		x"ffffffff", -- 1fb04
		x"ffffffff", -- 1fb08
		x"ffffffff", -- 1fb0c
		x"ffffffff", -- 1fb10
		x"ffffffff", -- 1fb14
		x"ffffffff", -- 1fb18
		x"ffffffff", -- 1fb1c
		x"ffffffff", -- 1fb20
		x"ffffffff", -- 1fb24
		x"ffffffff", -- 1fb28
		x"ffffffff", -- 1fb2c
		x"ffffffff", -- 1fb30
		x"ffffffff", -- 1fb34
		x"ffffffff", -- 1fb38
		x"ffffffff", -- 1fb3c
		x"ffffffff", -- 1fb40
		x"ffffffff", -- 1fb44
		x"ffffffff", -- 1fb48
		x"ffffffff", -- 1fb4c
		x"ffffffff", -- 1fb50
		x"ffffffff", -- 1fb54
		x"ffffffff", -- 1fb58
		x"ffffffff", -- 1fb5c
		x"ffffffff", -- 1fb60
		x"ffffffff", -- 1fb64
		x"ffffffff", -- 1fb68
		x"ffffffff", -- 1fb6c
		x"ffffffff", -- 1fb70
		x"ffffffff", -- 1fb74
		x"ffffffff", -- 1fb78
		x"ffffffff", -- 1fb7c
		x"ffffffff", -- 1fb80
		x"ffffffff", -- 1fb84
		x"ffffffff", -- 1fb88
		x"ffffffff", -- 1fb8c
		x"ffffffff", -- 1fb90
		x"ffffffff", -- 1fb94
		x"ffffffff", -- 1fb98
		x"ffffffff", -- 1fb9c
		x"ffffffff", -- 1fba0
		x"ffffffff", -- 1fba4
		x"ffffffff", -- 1fba8
		x"ffffffff", -- 1fbac
		x"ffffffff", -- 1fbb0
		x"ffffffff", -- 1fbb4
		x"ffffffff", -- 1fbb8
		x"ffffffff", -- 1fbbc
		x"ffffffff", -- 1fbc0
		x"ffffffff", -- 1fbc4
		x"ffffffff", -- 1fbc8
		x"ffffffff", -- 1fbcc
		x"ffffffff", -- 1fbd0
		x"ffffffff", -- 1fbd4
		x"ffffffff", -- 1fbd8
		x"ffffffff", -- 1fbdc
		x"ffffffff", -- 1fbe0
		x"ffffffff", -- 1fbe4
		x"ffffffff", -- 1fbe8
		x"ffffffff", -- 1fbec
		x"ffffffff", -- 1fbf0
		x"ffffffff", -- 1fbf4
		x"ffffffff", -- 1fbf8
		x"ffffffff", -- 1fbfc
		x"ffffffff", -- 1fc00
		x"ffffffff", -- 1fc04
		x"ffffffff", -- 1fc08
		x"ffffffff", -- 1fc0c
		x"ffffffff", -- 1fc10
		x"ffffffff", -- 1fc14
		x"ffffffff", -- 1fc18
		x"ffffffff", -- 1fc1c
		x"ffffffff", -- 1fc20
		x"ffffffff", -- 1fc24
		x"ffffffff", -- 1fc28
		x"ffffffff", -- 1fc2c
		x"ffffffff", -- 1fc30
		x"ffffffff", -- 1fc34
		x"ffffffff", -- 1fc38
		x"ffffffff", -- 1fc3c
		x"ffffffff", -- 1fc40
		x"ffffffff", -- 1fc44
		x"ffffffff", -- 1fc48
		x"ffffffff", -- 1fc4c
		x"ffffffff", -- 1fc50
		x"ffffffff", -- 1fc54
		x"ffffffff", -- 1fc58
		x"ffffffff", -- 1fc5c
		x"ffffffff", -- 1fc60
		x"ffffffff", -- 1fc64
		x"ffffffff", -- 1fc68
		x"ffffffff", -- 1fc6c
		x"ffffffff", -- 1fc70
		x"ffffffff", -- 1fc74
		x"ffffffff", -- 1fc78
		x"ffffffff", -- 1fc7c
		x"ffffffff", -- 1fc80
		x"ffffffff", -- 1fc84
		x"ffffffff", -- 1fc88
		x"ffffffff", -- 1fc8c
		x"ffffffff", -- 1fc90
		x"ffffffff", -- 1fc94
		x"ffffffff", -- 1fc98
		x"ffffffff", -- 1fc9c
		x"ffffffff", -- 1fca0
		x"ffffffff", -- 1fca4
		x"ffffffff", -- 1fca8
		x"ffffffff", -- 1fcac
		x"ffffffff", -- 1fcb0
		x"ffffffff", -- 1fcb4
		x"ffffffff", -- 1fcb8
		x"ffffffff", -- 1fcbc
		x"ffffffff", -- 1fcc0
		x"ffffffff", -- 1fcc4
		x"ffffffff", -- 1fcc8
		x"ffffffff", -- 1fccc
		x"ffffffff", -- 1fcd0
		x"ffffffff", -- 1fcd4
		x"ffffffff", -- 1fcd8
		x"ffffffff", -- 1fcdc
		x"ffffffff", -- 1fce0
		x"ffffffff", -- 1fce4
		x"ffffffff", -- 1fce8
		x"ffffffff", -- 1fcec
		x"ffffffff", -- 1fcf0
		x"ffffffff", -- 1fcf4
		x"ffffffff", -- 1fcf8
		x"ffffffff", -- 1fcfc
		x"ffffffff", -- 1fd00
		x"ffffffff", -- 1fd04
		x"ffffffff", -- 1fd08
		x"ffffffff", -- 1fd0c
		x"ffffffff", -- 1fd10
		x"ffffffff", -- 1fd14
		x"ffffffff", -- 1fd18
		x"ffffffff", -- 1fd1c
		x"ffffffff", -- 1fd20
		x"ffffffff", -- 1fd24
		x"ffffffff", -- 1fd28
		x"ffffffff", -- 1fd2c
		x"ffffffff", -- 1fd30
		x"ffffffff", -- 1fd34
		x"ffffffff", -- 1fd38
		x"ffffffff", -- 1fd3c
		x"ffffffff", -- 1fd40
		x"ffffffff", -- 1fd44
		x"ffffffff", -- 1fd48
		x"ffffffff", -- 1fd4c
		x"ffffffff", -- 1fd50
		x"ffffffff", -- 1fd54
		x"ffffffff", -- 1fd58
		x"ffffffff", -- 1fd5c
		x"ffffffff", -- 1fd60
		x"ffffffff", -- 1fd64
		x"ffffffff", -- 1fd68
		x"ffffffff", -- 1fd6c
		x"ffffffff", -- 1fd70
		x"ffffffff", -- 1fd74
		x"ffffffff", -- 1fd78
		x"ffffffff", -- 1fd7c
		x"ffffffff", -- 1fd80
		x"ffffffff", -- 1fd84
		x"ffffffff", -- 1fd88
		x"ffffffff", -- 1fd8c
		x"ffffffff", -- 1fd90
		x"ffffffff", -- 1fd94
		x"ffffffff", -- 1fd98
		x"ffffffff", -- 1fd9c
		x"ffffffff", -- 1fda0
		x"ffffffff", -- 1fda4
		x"ffffffff", -- 1fda8
		x"ffffffff", -- 1fdac
		x"ffffffff", -- 1fdb0
		x"ffffffff", -- 1fdb4
		x"ffffffff", -- 1fdb8
		x"ffffffff", -- 1fdbc
		x"ffffffff", -- 1fdc0
		x"ffffffff", -- 1fdc4
		x"ffffffff", -- 1fdc8
		x"ffffffff", -- 1fdcc
		x"ffffffff", -- 1fdd0
		x"ffffffff", -- 1fdd4
		x"ffffffff", -- 1fdd8
		x"ffffffff", -- 1fddc
		x"ffffffff", -- 1fde0
		x"ffffffff", -- 1fde4
		x"ffffffff", -- 1fde8
		x"ffffffff", -- 1fdec
		x"ffffffff", -- 1fdf0
		x"ffffffff", -- 1fdf4
		x"ffffffff", -- 1fdf8
		x"ffffffff", -- 1fdfc
		x"ffffffff", -- 1fe00
		x"ffffffff", -- 1fe04
		x"ffffffff", -- 1fe08
		x"ffffffff", -- 1fe0c
		x"ffffffff", -- 1fe10
		x"ffffffff", -- 1fe14
		x"ffffffff", -- 1fe18
		x"ffffffff", -- 1fe1c
		x"ffffffff", -- 1fe20
		x"ffffffff", -- 1fe24
		x"ffffffff", -- 1fe28
		x"ffffffff", -- 1fe2c
		x"ffffffff", -- 1fe30
		x"ffffffff", -- 1fe34
		x"ffffffff", -- 1fe38
		x"ffffffff", -- 1fe3c
		x"ffffffff", -- 1fe40
		x"ffffffff", -- 1fe44
		x"ffffffff", -- 1fe48
		x"ffffffff", -- 1fe4c
		x"ffffffff", -- 1fe50
		x"ffffffff", -- 1fe54
		x"ffffffff", -- 1fe58
		x"ffffffff", -- 1fe5c
		x"ffffffff", -- 1fe60
		x"ffffffff", -- 1fe64
		x"ffffffff", -- 1fe68
		x"ffffffff", -- 1fe6c
		x"ffffffff", -- 1fe70
		x"ffffffff", -- 1fe74
		x"ffffffff", -- 1fe78
		x"ffffffff", -- 1fe7c
		x"ffffffff", -- 1fe80
		x"ffffffff", -- 1fe84
		x"ffffffff", -- 1fe88
		x"ffffffff", -- 1fe8c
		x"ffffffff", -- 1fe90
		x"ffffffff", -- 1fe94
		x"ffffffff", -- 1fe98
		x"ffffffff", -- 1fe9c
		x"ffffffff", -- 1fea0
		x"ffffffff", -- 1fea4
		x"ffffffff", -- 1fea8
		x"ffffffff", -- 1feac
		x"ffffffff", -- 1feb0
		x"ffffffff", -- 1feb4
		x"ffffffff", -- 1feb8
		x"ffffffff", -- 1febc
		x"ffffffff", -- 1fec0
		x"ffffffff", -- 1fec4
		x"ffffffff", -- 1fec8
		x"ffffffff", -- 1fecc
		x"ffffffff", -- 1fed0
		x"ffffffff", -- 1fed4
		x"ffffffff", -- 1fed8
		x"ffffffff", -- 1fedc
		x"ffffffff", -- 1fee0
		x"ffffffff", -- 1fee4
		x"ffffffff", -- 1fee8
		x"ffffffff", -- 1feec
		x"ffffffff", -- 1fef0
		x"ffffffff", -- 1fef4
		x"ffffffff", -- 1fef8
		x"ffffffff", -- 1fefc
		x"ffffffff", -- 1ff00
		x"ffffffff", -- 1ff04
		x"ffffffff", -- 1ff08
		x"ffffffff", -- 1ff0c
		x"ffffffff", -- 1ff10
		x"ffffffff", -- 1ff14
		x"ffffffff", -- 1ff18
		x"ffffffff", -- 1ff1c
		x"ffffffff", -- 1ff20
		x"ffffffff", -- 1ff24
		x"ffffffff", -- 1ff28
		x"ffffffff", -- 1ff2c
		x"ffffffff", -- 1ff30
		x"ffffffff", -- 1ff34
		x"ffffffff", -- 1ff38
		x"ffffffff", -- 1ff3c
		x"ffffffff", -- 1ff40
		x"ffffffff", -- 1ff44
		x"ffffffff", -- 1ff48
		x"ffffffff", -- 1ff4c
		x"ffffffff", -- 1ff50
		x"ffffffff", -- 1ff54
		x"ffffffff", -- 1ff58
		x"ffffffff", -- 1ff5c
		x"ffffffff", -- 1ff60
		x"ffffffff", -- 1ff64
		x"ffffffff", -- 1ff68
		x"ffffffff", -- 1ff6c
		x"ffffffff", -- 1ff70
		x"ffffffff", -- 1ff74
		x"ffffffff", -- 1ff78
		x"ffffffff", -- 1ff7c
		x"ffffffff", -- 1ff80
		x"ffffffff", -- 1ff84
		x"ffffffff", -- 1ff88
		x"ffffffff", -- 1ff8c
		x"ffffffff", -- 1ff90
		x"ffffffff", -- 1ff94
		x"ffffffff", -- 1ff98
		x"ffffffff", -- 1ff9c
		x"ffffffff", -- 1ffa0
		x"ffffffff", -- 1ffa4
		x"ffffffff", -- 1ffa8
		x"ffffffff", -- 1ffac
		x"ffffffff", -- 1ffb0
		x"ffffffff", -- 1ffb4
		x"ffffffff", -- 1ffb8
		x"ffffffff", -- 1ffbc
		x"ffffffff", -- 1ffc0
		x"ffffffff", -- 1ffc4
		x"ffffffff", -- 1ffc8
		x"ffffffff", -- 1ffcc
		x"ffffffff", -- 1ffd0
		x"ffffffff", -- 1ffd4
		x"ffffffff", -- 1ffd8
		x"ffffffff", -- 1ffdc
		x"ffffffff", -- 1ffe0
		x"ffffffff", -- 1ffe4
		x"ffffffff", -- 1ffe8
		x"ffffffff", -- 1ffec
		x"ffffffff", -- 1fff0
		x"ffffffff", -- 1fff4
		x"ffffffff", -- 1fff8
		x"ffffffff"  -- 1fffc
);

begin
romp: process(clk_i)
begin
	if (rising_edge(clk_i)) then
		data_o <= rom_i(to_integer(unsigned(addr_i)));
	end if;
end process;
end rtl;
